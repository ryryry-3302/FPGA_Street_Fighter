module Gui_State1(
    input [12:0] pixel_index, 
    output reg [15:0] oled_colour 
); 

always@(pixel_index) 
begin
	case(pixel_index)
		0: oled_colour = 16'b00000_000000_00000;
		1: oled_colour = 16'b00000_000000_00000;
		2: oled_colour = 16'b00000_000000_00000;
		3: oled_colour = 16'b00000_000000_00000;
		4: oled_colour = 16'b00000_000000_00000;
		5: oled_colour = 16'b00000_000000_00000;
		6: oled_colour = 16'b00000_000000_00000;
		7: oled_colour = 16'b00000_000000_00000;
		8: oled_colour = 16'b00000_000000_00000;
		9: oled_colour = 16'b00000_000000_00000;
		10: oled_colour = 16'b00000_000000_00000;
		11: oled_colour = 16'b00000_000000_00000;
		12: oled_colour = 16'b00000_000000_00000;
		13: oled_colour = 16'b00000_000000_00000;
		14: oled_colour = 16'b00000_000000_00000;
		15: oled_colour = 16'b00000_000000_00000;
		16: oled_colour = 16'b00000_000000_00000;
		17: oled_colour = 16'b00000_000000_00000;
		18: oled_colour = 16'b00000_000000_00000;
		19: oled_colour = 16'b00000_000000_00000;
		20: oled_colour = 16'b00000_000000_00000;
		21: oled_colour = 16'b00000_000000_00000;
		22: oled_colour = 16'b00000_000000_00000;
		23: oled_colour = 16'b00000_000000_00000;
		24: oled_colour = 16'b00000_000000_00000;
		25: oled_colour = 16'b00000_000000_00000;
		26: oled_colour = 16'b00000_000000_00000;
		27: oled_colour = 16'b00000_000000_00000;
		28: oled_colour = 16'b00000_000000_00000;
		29: oled_colour = 16'b00000_000000_00000;
		30: oled_colour = 16'b00000_000000_00000;
		31: oled_colour = 16'b00000_000000_00000;
		32: oled_colour = 16'b00000_000000_00000;
		33: oled_colour = 16'b00000_000000_00000;
		34: oled_colour = 16'b00000_000000_00000;
		35: oled_colour = 16'b00000_000000_00000;
		36: oled_colour = 16'b00000_000000_00000;
		37: oled_colour = 16'b00000_000000_00000;
		38: oled_colour = 16'b00000_000000_00000;
		39: oled_colour = 16'b00000_000000_00000;
		40: oled_colour = 16'b00000_000000_00000;
		41: oled_colour = 16'b00000_000000_00000;
		42: oled_colour = 16'b00000_000000_00000;
		43: oled_colour = 16'b00000_000000_00000;
		44: oled_colour = 16'b00000_000000_00000;
		45: oled_colour = 16'b00000_000000_00000;
		46: oled_colour = 16'b00000_000000_00000;
		47: oled_colour = 16'b00000_000000_00000;
		48: oled_colour = 16'b00000_000000_00000;
		49: oled_colour = 16'b00000_000000_00000;
		50: oled_colour = 16'b00000_000000_00000;
		51: oled_colour = 16'b00000_000000_00000;
		52: oled_colour = 16'b00000_000000_00000;
		53: oled_colour = 16'b00000_000000_00000;
		54: oled_colour = 16'b00000_000000_00000;
		55: oled_colour = 16'b00000_000000_00000;
		56: oled_colour = 16'b00000_000000_00000;
		57: oled_colour = 16'b00000_000000_00000;
		58: oled_colour = 16'b00000_000000_00000;
		59: oled_colour = 16'b00000_000000_00000;
		60: oled_colour = 16'b00000_000000_00000;
		61: oled_colour = 16'b00000_000000_00000;
		62: oled_colour = 16'b00000_000000_00000;
		63: oled_colour = 16'b00000_000000_00000;
		64: oled_colour = 16'b00000_000000_00000;
		65: oled_colour = 16'b00000_000000_00000;
		66: oled_colour = 16'b00000_000000_00000;
		67: oled_colour = 16'b00000_000000_00000;
		68: oled_colour = 16'b00000_000000_00000;
		69: oled_colour = 16'b00000_000000_00000;
		70: oled_colour = 16'b00000_000000_00000;
		71: oled_colour = 16'b00000_000000_00000;
		72: oled_colour = 16'b00000_000000_00000;
		73: oled_colour = 16'b00000_000000_00000;
		74: oled_colour = 16'b00000_000000_00000;
		75: oled_colour = 16'b00000_000000_00000;
		76: oled_colour = 16'b00000_000000_00000;
		77: oled_colour = 16'b00000_000000_00000;
		78: oled_colour = 16'b00000_000000_00000;
		79: oled_colour = 16'b00000_000000_00000;
		80: oled_colour = 16'b00000_000000_00000;
		81: oled_colour = 16'b00000_000000_00000;
		82: oled_colour = 16'b00000_000000_00000;
		83: oled_colour = 16'b00000_000000_00000;
		84: oled_colour = 16'b00000_000000_00000;
		85: oled_colour = 16'b00000_000000_00000;
		86: oled_colour = 16'b00000_000000_00000;
		87: oled_colour = 16'b00000_000000_00000;
		88: oled_colour = 16'b00000_000000_00000;
		89: oled_colour = 16'b00000_000000_00000;
		90: oled_colour = 16'b00000_000000_00000;
		91: oled_colour = 16'b00000_000000_00000;
		92: oled_colour = 16'b00000_000000_00000;
		93: oled_colour = 16'b00000_000000_00000;
		94: oled_colour = 16'b00000_000000_00000;
		95: oled_colour = 16'b00000_000000_00000;
		96: oled_colour = 16'b00000_000000_00000;
		97: oled_colour = 16'b00000_000000_00000;
		98: oled_colour = 16'b00000_000000_00000;
		99: oled_colour = 16'b00000_000000_00000;
		100: oled_colour = 16'b00000_000000_00000;
		101: oled_colour = 16'b00000_000000_00000;
		102: oled_colour = 16'b00000_000000_00000;
		103: oled_colour = 16'b00000_000000_00000;
		104: oled_colour = 16'b00000_000000_00000;
		105: oled_colour = 16'b00000_000000_00000;
		106: oled_colour = 16'b00000_000000_00000;
		107: oled_colour = 16'b00000_000000_00000;
		108: oled_colour = 16'b00000_000000_00000;
		109: oled_colour = 16'b00000_000000_00000;
		110: oled_colour = 16'b00000_000000_00000;
		111: oled_colour = 16'b00000_000000_00000;
		112: oled_colour = 16'b00000_000000_00000;
		113: oled_colour = 16'b00000_000000_00000;
		114: oled_colour = 16'b00000_000000_00000;
		115: oled_colour = 16'b00000_000000_00000;
		116: oled_colour = 16'b00000_000000_00000;
		117: oled_colour = 16'b00000_000000_00000;
		118: oled_colour = 16'b00000_000000_00000;
		119: oled_colour = 16'b00000_000000_00000;
		120: oled_colour = 16'b00000_000000_00000;
		121: oled_colour = 16'b00000_000000_00000;
		122: oled_colour = 16'b00000_000000_00000;
		123: oled_colour = 16'b00000_000000_00000;
		124: oled_colour = 16'b00000_000000_00000;
		125: oled_colour = 16'b00000_000000_00000;
		126: oled_colour = 16'b00000_000000_00000;
		127: oled_colour = 16'b00000_000000_00000;
		128: oled_colour = 16'b00000_000000_00000;
		129: oled_colour = 16'b00000_000000_00000;
		130: oled_colour = 16'b00000_000000_00000;
		131: oled_colour = 16'b00000_000000_00000;
		132: oled_colour = 16'b00000_000000_00000;
		133: oled_colour = 16'b00000_000000_00000;
		134: oled_colour = 16'b00000_000000_00000;
		135: oled_colour = 16'b00000_000000_00000;
		136: oled_colour = 16'b00000_000000_00000;
		137: oled_colour = 16'b00000_000000_00000;
		138: oled_colour = 16'b00000_000000_00000;
		139: oled_colour = 16'b00000_000000_00000;
		140: oled_colour = 16'b00000_000000_00000;
		141: oled_colour = 16'b00000_000000_00000;
		142: oled_colour = 16'b00000_000000_00000;
		143: oled_colour = 16'b00000_000000_00000;
		144: oled_colour = 16'b00000_000000_00000;
		145: oled_colour = 16'b00000_000000_00000;
		146: oled_colour = 16'b00000_000000_00000;
		147: oled_colour = 16'b00000_000000_00000;
		148: oled_colour = 16'b00000_000000_00000;
		149: oled_colour = 16'b00000_000000_00000;
		150: oled_colour = 16'b00000_000000_00000;
		151: oled_colour = 16'b00000_000000_00000;
		152: oled_colour = 16'b00000_000000_00000;
		153: oled_colour = 16'b00000_000000_00000;
		154: oled_colour = 16'b00000_000000_00000;
		155: oled_colour = 16'b00000_000000_00000;
		156: oled_colour = 16'b00000_000000_00000;
		157: oled_colour = 16'b00000_000000_00000;
		158: oled_colour = 16'b00000_000000_00000;
		159: oled_colour = 16'b00000_000000_00000;
		160: oled_colour = 16'b00000_000000_00000;
		161: oled_colour = 16'b00000_000000_00000;
		162: oled_colour = 16'b00000_000000_00000;
		163: oled_colour = 16'b00000_000000_00000;
		164: oled_colour = 16'b00000_000000_00000;
		165: oled_colour = 16'b00000_000000_00000;
		166: oled_colour = 16'b00000_000000_00000;
		167: oled_colour = 16'b00000_000000_00000;
		168: oled_colour = 16'b00000_000000_00000;
		169: oled_colour = 16'b00000_000000_00000;
		170: oled_colour = 16'b00000_000000_00000;
		171: oled_colour = 16'b00000_000000_00000;
		172: oled_colour = 16'b00000_000000_00000;
		173: oled_colour = 16'b00000_000000_00000;
		174: oled_colour = 16'b00000_000000_00000;
		175: oled_colour = 16'b00000_000000_00000;
		176: oled_colour = 16'b00000_000000_00000;
		177: oled_colour = 16'b00000_000000_00000;
		178: oled_colour = 16'b00000_000000_00000;
		179: oled_colour = 16'b00000_000000_00000;
		180: oled_colour = 16'b00000_000000_00000;
		181: oled_colour = 16'b00000_000000_00000;
		182: oled_colour = 16'b00000_000000_00000;
		183: oled_colour = 16'b00000_000000_00000;
		184: oled_colour = 16'b00000_000000_00000;
		185: oled_colour = 16'b00000_000000_00000;
		186: oled_colour = 16'b00000_000000_00000;
		187: oled_colour = 16'b00000_000000_00000;
		188: oled_colour = 16'b00000_000000_00000;
		189: oled_colour = 16'b00000_000000_00000;
		190: oled_colour = 16'b00000_000000_00000;
		191: oled_colour = 16'b00000_000000_00000;
		192: oled_colour = 16'b00000_000000_00000;
		193: oled_colour = 16'b00000_000000_00000;
		194: oled_colour = 16'b00000_000000_00000;
		195: oled_colour = 16'b00000_000000_00000;
		196: oled_colour = 16'b00000_000000_00000;
		197: oled_colour = 16'b00000_000000_00000;
		198: oled_colour = 16'b00000_000000_00000;
		199: oled_colour = 16'b00000_000000_00000;
		200: oled_colour = 16'b00000_000000_00000;
		201: oled_colour = 16'b00000_000000_00000;
		202: oled_colour = 16'b00000_000000_00000;
		203: oled_colour = 16'b00000_000000_00000;
		204: oled_colour = 16'b00000_000000_00000;
		205: oled_colour = 16'b00000_000000_00000;
		206: oled_colour = 16'b00000_000000_00000;
		207: oled_colour = 16'b00000_000000_00000;
		208: oled_colour = 16'b00000_000000_00000;
		209: oled_colour = 16'b00000_000000_00000;
		210: oled_colour = 16'b00000_000000_00000;
		211: oled_colour = 16'b00000_000000_00000;
		212: oled_colour = 16'b00000_000000_00000;
		213: oled_colour = 16'b00000_000000_00000;
		214: oled_colour = 16'b00000_000000_00000;
		215: oled_colour = 16'b00000_000000_00000;
		216: oled_colour = 16'b00000_000000_00000;
		217: oled_colour = 16'b00000_000000_00000;
		218: oled_colour = 16'b00000_000000_00000;
		219: oled_colour = 16'b00000_000000_00000;
		220: oled_colour = 16'b00000_000000_00000;
		221: oled_colour = 16'b00000_000000_00000;
		222: oled_colour = 16'b00000_000000_00000;
		223: oled_colour = 16'b00000_000000_00000;
		224: oled_colour = 16'b00000_000000_00000;
		225: oled_colour = 16'b00000_000000_00000;
		226: oled_colour = 16'b00000_000000_00000;
		227: oled_colour = 16'b00000_000000_00000;
		228: oled_colour = 16'b00000_000000_00000;
		229: oled_colour = 16'b00000_000000_00000;
		230: oled_colour = 16'b00000_000000_00000;
		231: oled_colour = 16'b00000_000000_00000;
		232: oled_colour = 16'b00000_000000_00000;
		233: oled_colour = 16'b00000_000000_00000;
		234: oled_colour = 16'b00000_000000_00000;
		235: oled_colour = 16'b00000_000000_00000;
		236: oled_colour = 16'b00000_000000_00000;
		237: oled_colour = 16'b00000_000000_00000;
		238: oled_colour = 16'b00000_000000_00000;
		239: oled_colour = 16'b00000_000000_00000;
		240: oled_colour = 16'b00000_000000_00000;
		241: oled_colour = 16'b00000_000000_00000;
		242: oled_colour = 16'b00000_000000_00000;
		243: oled_colour = 16'b00000_000000_00000;
		244: oled_colour = 16'b00000_000000_00000;
		245: oled_colour = 16'b00000_000000_00000;
		246: oled_colour = 16'b00000_000000_00000;
		247: oled_colour = 16'b00000_000000_00000;
		248: oled_colour = 16'b00000_000000_00000;
		249: oled_colour = 16'b00000_000000_00000;
		250: oled_colour = 16'b00000_000000_00000;
		251: oled_colour = 16'b00000_000000_00000;
		252: oled_colour = 16'b00000_000000_00000;
		253: oled_colour = 16'b00000_000000_00000;
		254: oled_colour = 16'b00000_000000_00000;
		255: oled_colour = 16'b00000_000000_00000;
		256: oled_colour = 16'b00000_000000_00000;
		257: oled_colour = 16'b00000_000000_00000;
		258: oled_colour = 16'b00000_000000_00000;
		259: oled_colour = 16'b00000_000000_00000;
		260: oled_colour = 16'b00000_000000_00000;
		261: oled_colour = 16'b00000_000000_00000;
		262: oled_colour = 16'b00000_000000_00000;
		263: oled_colour = 16'b00000_000000_00000;
		264: oled_colour = 16'b00000_000000_00000;
		265: oled_colour = 16'b00000_000000_00000;
		266: oled_colour = 16'b00000_000000_00000;
		267: oled_colour = 16'b00000_000000_00000;
		268: oled_colour = 16'b00000_000000_00000;
		269: oled_colour = 16'b00000_000000_00000;
		270: oled_colour = 16'b00000_000000_00000;
		271: oled_colour = 16'b00000_000000_00000;
		272: oled_colour = 16'b00000_000000_00000;
		273: oled_colour = 16'b00000_000000_00000;
		274: oled_colour = 16'b00000_000000_00000;
		275: oled_colour = 16'b00000_000000_00000;
		276: oled_colour = 16'b00000_000000_00000;
		277: oled_colour = 16'b00000_000000_00000;
		278: oled_colour = 16'b00000_000000_00000;
		279: oled_colour = 16'b00000_000000_00000;
		280: oled_colour = 16'b00000_000000_00000;
		281: oled_colour = 16'b00000_000000_00000;
		282: oled_colour = 16'b00000_000000_00000;
		283: oled_colour = 16'b00000_000000_00000;
		284: oled_colour = 16'b00000_000000_00000;
		285: oled_colour = 16'b00000_000000_00000;
		286: oled_colour = 16'b00000_000000_00000;
		287: oled_colour = 16'b00000_000000_00000;
		288: oled_colour = 16'b00000_000000_00000;
		289: oled_colour = 16'b00000_000000_00000;
		290: oled_colour = 16'b00000_000000_00000;
		291: oled_colour = 16'b00000_000000_00000;
		292: oled_colour = 16'b00000_000000_00000;
		293: oled_colour = 16'b00000_000000_00000;
		294: oled_colour = 16'b00000_000000_00000;
		295: oled_colour = 16'b00000_000000_00000;
		296: oled_colour = 16'b00000_000000_00000;
		297: oled_colour = 16'b00000_000000_00000;
		298: oled_colour = 16'b00000_000000_00000;
		299: oled_colour = 16'b00000_000000_00000;
		300: oled_colour = 16'b00000_000000_00000;
		301: oled_colour = 16'b00000_000000_00000;
		302: oled_colour = 16'b00000_000000_00000;
		303: oled_colour = 16'b00000_000000_00000;
		304: oled_colour = 16'b00000_000000_00000;
		305: oled_colour = 16'b00000_000000_00000;
		306: oled_colour = 16'b00000_000000_00000;
		307: oled_colour = 16'b00000_000000_00000;
		308: oled_colour = 16'b00000_000000_00000;
		309: oled_colour = 16'b00000_000000_00000;
		310: oled_colour = 16'b00000_000000_00000;
		311: oled_colour = 16'b00000_000000_00000;
		312: oled_colour = 16'b00000_000000_00000;
		313: oled_colour = 16'b00000_000000_00000;
		314: oled_colour = 16'b00000_000000_00000;
		315: oled_colour = 16'b00000_000000_00000;
		316: oled_colour = 16'b00000_000000_00000;
		317: oled_colour = 16'b00000_000000_00000;
		318: oled_colour = 16'b00000_000000_00000;
		319: oled_colour = 16'b00000_000000_00000;
		320: oled_colour = 16'b00000_000000_00000;
		321: oled_colour = 16'b00000_000000_00000;
		322: oled_colour = 16'b00000_000000_00000;
		323: oled_colour = 16'b00000_000000_00000;
		324: oled_colour = 16'b00000_000000_00000;
		325: oled_colour = 16'b00000_000000_00000;
		326: oled_colour = 16'b00000_000000_00000;
		327: oled_colour = 16'b00000_000000_00000;
		328: oled_colour = 16'b00000_000000_00000;
		329: oled_colour = 16'b00000_000000_00000;
		330: oled_colour = 16'b00000_000000_00000;
		331: oled_colour = 16'b00000_000000_00000;
		332: oled_colour = 16'b00000_000000_00000;
		333: oled_colour = 16'b00000_000000_00000;
		334: oled_colour = 16'b00000_000000_00000;
		335: oled_colour = 16'b00000_000000_00000;
		336: oled_colour = 16'b00000_000000_00000;
		337: oled_colour = 16'b00000_000000_00000;
		338: oled_colour = 16'b00000_000000_00000;
		339: oled_colour = 16'b00000_000000_00000;
		340: oled_colour = 16'b00000_000000_00000;
		341: oled_colour = 16'b00000_000000_00000;
		342: oled_colour = 16'b00000_000000_00000;
		343: oled_colour = 16'b00000_000000_00000;
		344: oled_colour = 16'b00000_000000_00000;
		345: oled_colour = 16'b00000_000000_00000;
		346: oled_colour = 16'b00000_000000_00000;
		347: oled_colour = 16'b00000_000000_00000;
		348: oled_colour = 16'b00000_000000_00000;
		349: oled_colour = 16'b00000_000000_00000;
		350: oled_colour = 16'b00000_000000_00000;
		351: oled_colour = 16'b00000_000000_00000;
		352: oled_colour = 16'b00000_000000_00000;
		353: oled_colour = 16'b00000_000000_00000;
		354: oled_colour = 16'b00000_000000_00000;
		355: oled_colour = 16'b00000_000000_00000;
		356: oled_colour = 16'b00000_000000_00000;
		357: oled_colour = 16'b00000_000000_00000;
		358: oled_colour = 16'b00000_000000_00000;
		359: oled_colour = 16'b00000_000000_00000;
		360: oled_colour = 16'b00000_000000_00000;
		361: oled_colour = 16'b00000_000000_00000;
		362: oled_colour = 16'b00000_000000_00000;
		363: oled_colour = 16'b00000_000000_00000;
		364: oled_colour = 16'b00000_000000_00000;
		365: oled_colour = 16'b00000_000000_00000;
		366: oled_colour = 16'b00000_000000_00000;
		367: oled_colour = 16'b00000_000000_00000;
		368: oled_colour = 16'b00000_000000_00000;
		369: oled_colour = 16'b00000_000000_00000;
		370: oled_colour = 16'b00000_000000_00000;
		371: oled_colour = 16'b00000_000000_00000;
		372: oled_colour = 16'b00000_000000_00000;
		373: oled_colour = 16'b00000_000000_00000;
		374: oled_colour = 16'b00000_000000_00000;
		375: oled_colour = 16'b00000_000000_00000;
		376: oled_colour = 16'b00000_000000_00000;
		377: oled_colour = 16'b00000_000000_00000;
		378: oled_colour = 16'b00000_000000_00000;
		379: oled_colour = 16'b00000_000000_00000;
		380: oled_colour = 16'b00000_000000_00000;
		381: oled_colour = 16'b00000_000000_00000;
		382: oled_colour = 16'b00000_000000_00000;
		383: oled_colour = 16'b00000_000000_00000;
		384: oled_colour = 16'b00000_000000_00000;
		385: oled_colour = 16'b00000_000000_00000;
		386: oled_colour = 16'b00000_000000_00000;
		387: oled_colour = 16'b00000_000000_00000;
		388: oled_colour = 16'b00000_000000_00000;
		389: oled_colour = 16'b00000_000000_00000;
		390: oled_colour = 16'b00000_000000_00000;
		391: oled_colour = 16'b00000_000000_00000;
		392: oled_colour = 16'b00000_000000_00000;
		393: oled_colour = 16'b00000_000000_00000;
		394: oled_colour = 16'b00000_000000_00000;
		395: oled_colour = 16'b00000_000000_00000;
		396: oled_colour = 16'b00000_000000_00000;
		397: oled_colour = 16'b00000_000000_00000;
		398: oled_colour = 16'b00000_000000_00000;
		399: oled_colour = 16'b00000_000000_00000;
		400: oled_colour = 16'b00000_000000_00000;
		401: oled_colour = 16'b00000_000000_00000;
		402: oled_colour = 16'b00000_000000_00000;
		403: oled_colour = 16'b00000_000000_00000;
		404: oled_colour = 16'b00000_000000_00000;
		405: oled_colour = 16'b00000_000000_00000;
		406: oled_colour = 16'b00000_000000_00000;
		407: oled_colour = 16'b00000_000000_00000;
		408: oled_colour = 16'b00000_000000_00000;
		409: oled_colour = 16'b00000_000000_00000;
		410: oled_colour = 16'b00000_000000_00000;
		411: oled_colour = 16'b00000_000000_00000;
		412: oled_colour = 16'b00000_000000_00000;
		413: oled_colour = 16'b00000_000000_00000;
		414: oled_colour = 16'b00000_000000_00000;
		415: oled_colour = 16'b00000_000000_00000;
		416: oled_colour = 16'b00000_000000_00000;
		417: oled_colour = 16'b00000_000000_00000;
		418: oled_colour = 16'b00000_000000_00000;
		419: oled_colour = 16'b00000_000000_00000;
		420: oled_colour = 16'b00000_000000_00000;
		421: oled_colour = 16'b00000_000000_00000;
		422: oled_colour = 16'b00000_000000_00000;
		423: oled_colour = 16'b00000_000000_00000;
		424: oled_colour = 16'b00000_000000_00000;
		425: oled_colour = 16'b00000_000000_00000;
		426: oled_colour = 16'b00000_000000_00000;
		427: oled_colour = 16'b00000_000000_00000;
		428: oled_colour = 16'b00000_000000_00000;
		429: oled_colour = 16'b00000_000000_00000;
		430: oled_colour = 16'b00000_000000_00000;
		431: oled_colour = 16'b00000_000000_00000;
		432: oled_colour = 16'b00000_000000_00000;
		433: oled_colour = 16'b00000_000000_00000;
		434: oled_colour = 16'b00000_000000_00000;
		435: oled_colour = 16'b00000_000000_00000;
		436: oled_colour = 16'b00000_000000_00000;
		437: oled_colour = 16'b00000_000000_00000;
		438: oled_colour = 16'b00000_000000_00000;
		439: oled_colour = 16'b00000_000000_00000;
		440: oled_colour = 16'b00000_000000_00000;
		441: oled_colour = 16'b00000_000000_00000;
		442: oled_colour = 16'b00000_000000_00000;
		443: oled_colour = 16'b00000_000000_00000;
		444: oled_colour = 16'b00000_000000_00000;
		445: oled_colour = 16'b00000_000000_00000;
		446: oled_colour = 16'b00000_000000_00000;
		447: oled_colour = 16'b00000_000000_00000;
		448: oled_colour = 16'b00000_000000_00000;
		449: oled_colour = 16'b00000_000000_00000;
		450: oled_colour = 16'b00000_000000_00000;
		451: oled_colour = 16'b00000_000000_00000;
		452: oled_colour = 16'b00000_000000_00000;
		453: oled_colour = 16'b00000_000000_00000;
		454: oled_colour = 16'b00000_000000_00000;
		455: oled_colour = 16'b00000_000000_00000;
		456: oled_colour = 16'b00000_000000_00000;
		457: oled_colour = 16'b00000_000000_00000;
		458: oled_colour = 16'b00000_000000_00000;
		459: oled_colour = 16'b00000_000000_00000;
		460: oled_colour = 16'b00000_000000_00000;
		461: oled_colour = 16'b00000_000000_00000;
		462: oled_colour = 16'b00000_000000_00000;
		463: oled_colour = 16'b00000_000000_00000;
		464: oled_colour = 16'b00000_000000_00000;
		465: oled_colour = 16'b00000_000000_00000;
		466: oled_colour = 16'b00000_000000_00000;
		467: oled_colour = 16'b00000_000000_00000;
		468: oled_colour = 16'b00000_000000_00000;
		469: oled_colour = 16'b00000_000000_00000;
		470: oled_colour = 16'b00000_000000_00000;
		471: oled_colour = 16'b00000_000000_00000;
		472: oled_colour = 16'b00000_000000_00000;
		473: oled_colour = 16'b00000_000000_00000;
		474: oled_colour = 16'b00000_000000_00000;
		475: oled_colour = 16'b00000_000000_00000;
		476: oled_colour = 16'b00000_000000_00000;
		477: oled_colour = 16'b00000_000000_00000;
		478: oled_colour = 16'b00000_000000_00000;
		479: oled_colour = 16'b00000_000000_00000;
		480: oled_colour = 16'b00000_000000_00000;
		481: oled_colour = 16'b00000_000000_00000;
		482: oled_colour = 16'b00000_000000_00000;
		483: oled_colour = 16'b00000_000000_00000;
		484: oled_colour = 16'b00000_000000_00000;
		485: oled_colour = 16'b00000_000000_00000;
		486: oled_colour = 16'b00000_000000_00000;
		487: oled_colour = 16'b00000_000000_00000;
		488: oled_colour = 16'b00000_000000_00000;
		489: oled_colour = 16'b00000_000000_00000;
		490: oled_colour = 16'b00000_000000_00000;
		491: oled_colour = 16'b00000_000000_00000;
		492: oled_colour = 16'b00000_000000_00000;
		493: oled_colour = 16'b00000_000000_00000;
		494: oled_colour = 16'b00000_000000_00000;
		495: oled_colour = 16'b00000_000000_00000;
		496: oled_colour = 16'b00000_000000_00000;
		497: oled_colour = 16'b00000_000000_00000;
		498: oled_colour = 16'b00000_000000_00000;
		499: oled_colour = 16'b00000_000000_00000;
		500: oled_colour = 16'b00000_000000_00000;
		501: oled_colour = 16'b00000_000000_00000;
		502: oled_colour = 16'b00000_000000_00000;
		503: oled_colour = 16'b00000_000000_00000;
		504: oled_colour = 16'b00000_000000_00000;
		505: oled_colour = 16'b00000_000000_00000;
		506: oled_colour = 16'b00000_000000_00000;
		507: oled_colour = 16'b00000_000000_00000;
		508: oled_colour = 16'b00000_000000_00000;
		509: oled_colour = 16'b00000_000000_00000;
		510: oled_colour = 16'b00000_000000_00000;
		511: oled_colour = 16'b00000_000000_00000;
		512: oled_colour = 16'b00000_000000_00000;
		513: oled_colour = 16'b00000_000000_00000;
		514: oled_colour = 16'b00000_000000_00000;
		515: oled_colour = 16'b00000_000000_00000;
		516: oled_colour = 16'b00000_000000_00000;
		517: oled_colour = 16'b00000_000000_00000;
		518: oled_colour = 16'b00000_000000_00000;
		519: oled_colour = 16'b00000_000000_00000;
		520: oled_colour = 16'b00000_000000_00000;
		521: oled_colour = 16'b00000_000000_00000;
		522: oled_colour = 16'b00000_000000_00000;
		523: oled_colour = 16'b00000_000000_00000;
		524: oled_colour = 16'b00000_000000_00000;
		525: oled_colour = 16'b00000_000000_00000;
		526: oled_colour = 16'b00000_000000_00000;
		527: oled_colour = 16'b00000_000000_00000;
		528: oled_colour = 16'b00000_000000_00000;
		529: oled_colour = 16'b00000_000000_00000;
		530: oled_colour = 16'b00000_000000_00000;
		531: oled_colour = 16'b00000_000000_00000;
		532: oled_colour = 16'b00000_000000_00000;
		533: oled_colour = 16'b00000_000000_00000;
		534: oled_colour = 16'b00000_000000_00000;
		535: oled_colour = 16'b00000_000000_00000;
		536: oled_colour = 16'b00000_000000_00000;
		537: oled_colour = 16'b00000_000000_00000;
		538: oled_colour = 16'b00000_000000_00000;
		539: oled_colour = 16'b00000_000000_00000;
		540: oled_colour = 16'b00000_000000_00000;
		541: oled_colour = 16'b00000_000000_00000;
		542: oled_colour = 16'b00000_000000_00000;
		543: oled_colour = 16'b00000_000000_00000;
		544: oled_colour = 16'b00000_000000_00000;
		545: oled_colour = 16'b00000_000000_00000;
		546: oled_colour = 16'b00000_000000_00000;
		547: oled_colour = 16'b00000_000000_00000;
		548: oled_colour = 16'b00000_000000_00000;
		549: oled_colour = 16'b00000_000000_00000;
		550: oled_colour = 16'b00000_000000_00000;
		551: oled_colour = 16'b00000_000000_00000;
		552: oled_colour = 16'b00000_000000_00000;
		553: oled_colour = 16'b00000_000000_00000;
		554: oled_colour = 16'b00000_000000_00000;
		555: oled_colour = 16'b00000_000000_00000;
		556: oled_colour = 16'b00000_000000_00000;
		557: oled_colour = 16'b00000_000000_00000;
		558: oled_colour = 16'b00000_000000_00000;
		559: oled_colour = 16'b00000_000000_00000;
		560: oled_colour = 16'b00000_000000_00000;
		561: oled_colour = 16'b00000_000000_00000;
		562: oled_colour = 16'b00000_000000_00000;
		563: oled_colour = 16'b00000_000000_00000;
		564: oled_colour = 16'b00000_000000_00000;
		565: oled_colour = 16'b00000_000000_00000;
		566: oled_colour = 16'b00000_000000_00000;
		567: oled_colour = 16'b00000_000000_00000;
		568: oled_colour = 16'b00000_000000_00000;
		569: oled_colour = 16'b00000_000000_00000;
		570: oled_colour = 16'b00000_000000_00000;
		571: oled_colour = 16'b00000_000000_00000;
		572: oled_colour = 16'b00000_000000_00000;
		573: oled_colour = 16'b00000_000000_00000;
		574: oled_colour = 16'b00000_000000_00000;
		575: oled_colour = 16'b00000_000000_00000;
		576: oled_colour = 16'b00000_000000_00000;
		577: oled_colour = 16'b00000_000000_00000;
		578: oled_colour = 16'b00000_000000_00000;
		579: oled_colour = 16'b00000_000000_00000;
		580: oled_colour = 16'b00000_000000_00000;
		581: oled_colour = 16'b00000_000000_00000;
		582: oled_colour = 16'b00000_000000_00000;
		583: oled_colour = 16'b00000_000000_00000;
		584: oled_colour = 16'b00000_000000_00000;
		585: oled_colour = 16'b00000_000000_00000;
		586: oled_colour = 16'b00000_000000_00000;
		587: oled_colour = 16'b00000_000000_00000;
		588: oled_colour = 16'b00000_000000_00000;
		589: oled_colour = 16'b00000_000000_00000;
		590: oled_colour = 16'b00000_000000_00000;
		591: oled_colour = 16'b00000_000000_00000;
		592: oled_colour = 16'b00000_000000_00000;
		593: oled_colour = 16'b00000_000000_00000;
		594: oled_colour = 16'b00000_000000_00000;
		595: oled_colour = 16'b00000_000000_00000;
		596: oled_colour = 16'b00000_000000_00000;
		597: oled_colour = 16'b00000_000000_00000;
		598: oled_colour = 16'b00000_000000_00000;
		599: oled_colour = 16'b00000_000000_00000;
		600: oled_colour = 16'b00000_000000_00000;
		601: oled_colour = 16'b00000_000000_00000;
		602: oled_colour = 16'b00000_000000_00000;
		603: oled_colour = 16'b00000_000000_00000;
		604: oled_colour = 16'b00000_000000_00000;
		605: oled_colour = 16'b00000_000000_00000;
		606: oled_colour = 16'b00000_000000_00000;
		607: oled_colour = 16'b00000_000000_00000;
		608: oled_colour = 16'b00000_000000_00000;
		609: oled_colour = 16'b00000_000000_00000;
		610: oled_colour = 16'b00000_000000_00000;
		611: oled_colour = 16'b00000_000000_00000;
		612: oled_colour = 16'b00000_000000_00000;
		613: oled_colour = 16'b00000_000000_00000;
		614: oled_colour = 16'b00000_000000_00000;
		615: oled_colour = 16'b00000_000000_00000;
		616: oled_colour = 16'b00000_000000_00000;
		617: oled_colour = 16'b00000_000000_00000;
		618: oled_colour = 16'b00000_000000_00000;
		619: oled_colour = 16'b00000_000000_00000;
		620: oled_colour = 16'b00000_000000_00000;
		621: oled_colour = 16'b00000_000000_00000;
		622: oled_colour = 16'b00000_000000_00000;
		623: oled_colour = 16'b00000_000000_00000;
		624: oled_colour = 16'b00000_000000_00000;
		625: oled_colour = 16'b00000_000000_00000;
		626: oled_colour = 16'b00000_000000_00000;
		627: oled_colour = 16'b00000_000000_00000;
		628: oled_colour = 16'b00000_000000_00000;
		629: oled_colour = 16'b00000_000000_00000;
		630: oled_colour = 16'b00000_000000_00000;
		631: oled_colour = 16'b00000_000000_00000;
		632: oled_colour = 16'b00000_000000_00000;
		633: oled_colour = 16'b00000_000000_00000;
		634: oled_colour = 16'b00000_000000_00000;
		635: oled_colour = 16'b00000_000000_00000;
		636: oled_colour = 16'b00000_000000_00000;
		637: oled_colour = 16'b00000_000000_00000;
		638: oled_colour = 16'b00000_000000_00000;
		639: oled_colour = 16'b00000_000000_00000;
		640: oled_colour = 16'b00000_000000_00000;
		641: oled_colour = 16'b00000_000000_00000;
		642: oled_colour = 16'b00000_000000_00000;
		643: oled_colour = 16'b00000_000000_00000;
		644: oled_colour = 16'b00000_000000_00000;
		645: oled_colour = 16'b00000_000000_00000;
		646: oled_colour = 16'b00000_000000_00000;
		647: oled_colour = 16'b00000_000000_00000;
		648: oled_colour = 16'b00000_000000_00000;
		649: oled_colour = 16'b00000_000000_00000;
		650: oled_colour = 16'b00000_000000_00000;
		651: oled_colour = 16'b00000_000000_00000;
		652: oled_colour = 16'b00000_000000_00000;
		653: oled_colour = 16'b00000_000000_00000;
		654: oled_colour = 16'b00000_000000_00000;
		655: oled_colour = 16'b00000_000000_00000;
		656: oled_colour = 16'b00000_000000_00000;
		657: oled_colour = 16'b00000_000000_00000;
		658: oled_colour = 16'b00000_000000_00000;
		659: oled_colour = 16'b00000_000000_00000;
		660: oled_colour = 16'b00000_000000_00000;
		661: oled_colour = 16'b00000_000000_00000;
		662: oled_colour = 16'b00000_000000_00000;
		663: oled_colour = 16'b00000_000000_00000;
		664: oled_colour = 16'b00000_000000_00000;
		665: oled_colour = 16'b00000_000000_00000;
		666: oled_colour = 16'b00000_000000_00000;
		667: oled_colour = 16'b00000_000000_00000;
		668: oled_colour = 16'b00000_000000_00000;
		669: oled_colour = 16'b00000_000000_00000;
		670: oled_colour = 16'b00000_000000_00000;
		671: oled_colour = 16'b00000_000000_00000;
		672: oled_colour = 16'b00000_000000_00000;
		673: oled_colour = 16'b00000_000000_00000;
		674: oled_colour = 16'b00000_000000_00000;
		675: oled_colour = 16'b00000_000000_00000;
		676: oled_colour = 16'b00000_000000_00000;
		677: oled_colour = 16'b00000_000000_00000;
		678: oled_colour = 16'b00000_000000_00000;
		679: oled_colour = 16'b00000_000000_00000;
		680: oled_colour = 16'b00000_000000_00000;
		681: oled_colour = 16'b00000_000000_00000;
		682: oled_colour = 16'b00000_000000_00000;
		683: oled_colour = 16'b00000_000000_00000;
		684: oled_colour = 16'b00000_000000_00000;
		685: oled_colour = 16'b00000_000000_00000;
		686: oled_colour = 16'b00000_000000_00000;
		687: oled_colour = 16'b00000_000000_00000;
		688: oled_colour = 16'b00000_000000_00000;
		689: oled_colour = 16'b00000_000000_00000;
		690: oled_colour = 16'b00000_000000_00000;
		691: oled_colour = 16'b00000_000000_00000;
		692: oled_colour = 16'b00000_000000_00000;
		693: oled_colour = 16'b00000_000000_00000;
		694: oled_colour = 16'b00000_000000_00000;
		695: oled_colour = 16'b00000_000000_00000;
		696: oled_colour = 16'b00000_000000_00000;
		697: oled_colour = 16'b00000_000000_00000;
		698: oled_colour = 16'b00000_000000_00000;
		699: oled_colour = 16'b00000_000000_00000;
		700: oled_colour = 16'b00000_000000_00000;
		701: oled_colour = 16'b00000_000000_00000;
		702: oled_colour = 16'b00000_000000_00000;
		703: oled_colour = 16'b00000_000000_00000;
		704: oled_colour = 16'b00000_000000_00000;
		705: oled_colour = 16'b00000_000000_00000;
		706: oled_colour = 16'b00000_000000_00000;
		707: oled_colour = 16'b00000_000000_00000;
		708: oled_colour = 16'b00000_000000_00000;
		709: oled_colour = 16'b00000_000000_00000;
		710: oled_colour = 16'b00000_000000_00000;
		711: oled_colour = 16'b00000_000000_00000;
		712: oled_colour = 16'b00000_000000_00000;
		713: oled_colour = 16'b00000_000000_00000;
		714: oled_colour = 16'b00000_000000_00000;
		715: oled_colour = 16'b00000_000000_00000;
		716: oled_colour = 16'b00000_000000_00000;
		717: oled_colour = 16'b00000_000000_00000;
		718: oled_colour = 16'b00000_000000_00000;
		719: oled_colour = 16'b00000_000000_00000;
		720: oled_colour = 16'b00000_000000_00000;
		721: oled_colour = 16'b00000_000000_00000;
		722: oled_colour = 16'b00000_000000_00000;
		723: oled_colour = 16'b00000_000000_00000;
		724: oled_colour = 16'b00000_000000_00000;
		725: oled_colour = 16'b00000_000000_00000;
		726: oled_colour = 16'b00000_000000_00000;
		727: oled_colour = 16'b00000_000000_00000;
		728: oled_colour = 16'b00000_000000_00000;
		729: oled_colour = 16'b00000_000000_00000;
		730: oled_colour = 16'b00000_000000_00000;
		731: oled_colour = 16'b00000_000000_00000;
		732: oled_colour = 16'b00000_000000_00000;
		733: oled_colour = 16'b00000_000000_00000;
		734: oled_colour = 16'b00000_000000_00000;
		735: oled_colour = 16'b00000_000000_00000;
		736: oled_colour = 16'b00000_000000_00000;
		737: oled_colour = 16'b00000_000000_00000;
		738: oled_colour = 16'b00000_000000_00000;
		739: oled_colour = 16'b00000_000000_00000;
		740: oled_colour = 16'b00000_000000_00000;
		741: oled_colour = 16'b00000_000000_00000;
		742: oled_colour = 16'b00000_000000_00000;
		743: oled_colour = 16'b00000_000000_00000;
		744: oled_colour = 16'b00000_000000_00000;
		745: oled_colour = 16'b00000_000000_00000;
		746: oled_colour = 16'b00000_000000_00000;
		747: oled_colour = 16'b00000_000000_00000;
		748: oled_colour = 16'b00000_000000_00000;
		749: oled_colour = 16'b00000_000000_00000;
		750: oled_colour = 16'b00000_000000_00000;
		751: oled_colour = 16'b00000_000000_00000;
		752: oled_colour = 16'b00000_000000_00000;
		753: oled_colour = 16'b00000_000000_00000;
		754: oled_colour = 16'b00000_000000_00000;
		755: oled_colour = 16'b00000_000000_00000;
		756: oled_colour = 16'b00000_000000_00000;
		757: oled_colour = 16'b00000_000000_00000;
		758: oled_colour = 16'b00000_000000_00000;
		759: oled_colour = 16'b00000_000000_00000;
		760: oled_colour = 16'b00000_000000_00000;
		761: oled_colour = 16'b00000_000000_00000;
		762: oled_colour = 16'b00000_000000_00000;
		763: oled_colour = 16'b00000_000000_00000;
		764: oled_colour = 16'b00000_000000_00000;
		765: oled_colour = 16'b00000_000000_00000;
		766: oled_colour = 16'b00000_000000_00000;
		767: oled_colour = 16'b00000_000000_00000;
		768: oled_colour = 16'b00000_000000_00000;
		769: oled_colour = 16'b00000_000000_00000;
		770: oled_colour = 16'b00000_000000_00000;
		771: oled_colour = 16'b00000_000000_00000;
		772: oled_colour = 16'b00000_000000_00000;
		773: oled_colour = 16'b00000_000000_00000;
		774: oled_colour = 16'b00000_000000_00000;
		775: oled_colour = 16'b00000_000000_00000;
		776: oled_colour = 16'b00000_000000_00000;
		777: oled_colour = 16'b00000_000000_00000;
		778: oled_colour = 16'b00000_000000_00000;
		779: oled_colour = 16'b00000_000000_00000;
		780: oled_colour = 16'b00000_000000_00000;
		781: oled_colour = 16'b00000_000000_00000;
		782: oled_colour = 16'b00000_000000_00000;
		783: oled_colour = 16'b00000_000000_00000;
		784: oled_colour = 16'b00000_000000_00000;
		785: oled_colour = 16'b00000_000000_00000;
		786: oled_colour = 16'b00000_000000_00000;
		787: oled_colour = 16'b00000_000000_00000;
		788: oled_colour = 16'b00000_000000_00000;
		789: oled_colour = 16'b00000_000000_00000;
		790: oled_colour = 16'b00000_000000_00000;
		791: oled_colour = 16'b00000_000000_00000;
		792: oled_colour = 16'b00000_000000_00000;
		793: oled_colour = 16'b00000_000000_00000;
		794: oled_colour = 16'b00000_000000_00000;
		795: oled_colour = 16'b00000_000000_00000;
		796: oled_colour = 16'b00000_000000_00000;
		797: oled_colour = 16'b00000_000000_00000;
		798: oled_colour = 16'b00000_000000_00000;
		799: oled_colour = 16'b00000_000000_00000;
		800: oled_colour = 16'b00000_000000_00000;
		801: oled_colour = 16'b00000_000000_00000;
		802: oled_colour = 16'b00000_000000_00000;
		803: oled_colour = 16'b00000_000000_00000;
		804: oled_colour = 16'b00000_000000_00000;
		805: oled_colour = 16'b00000_000000_00000;
		806: oled_colour = 16'b00000_000000_00000;
		807: oled_colour = 16'b00000_000000_00000;
		808: oled_colour = 16'b00000_000000_00000;
		809: oled_colour = 16'b00000_000000_00000;
		810: oled_colour = 16'b00000_000000_00000;
		811: oled_colour = 16'b00000_000000_00000;
		812: oled_colour = 16'b00000_000000_00000;
		813: oled_colour = 16'b00000_000000_00000;
		814: oled_colour = 16'b00000_000000_00000;
		815: oled_colour = 16'b00000_000000_00000;
		816: oled_colour = 16'b00000_000000_00000;
		817: oled_colour = 16'b00000_000000_00000;
		818: oled_colour = 16'b00000_000000_00000;
		819: oled_colour = 16'b00000_000000_00000;
		820: oled_colour = 16'b00000_000000_00000;
		821: oled_colour = 16'b00000_000000_00000;
		822: oled_colour = 16'b00000_000000_00000;
		823: oled_colour = 16'b00000_000000_00000;
		824: oled_colour = 16'b00000_000000_00000;
		825: oled_colour = 16'b00000_000000_00000;
		826: oled_colour = 16'b00000_000000_00000;
		827: oled_colour = 16'b00000_000000_00000;
		828: oled_colour = 16'b00000_000000_00000;
		829: oled_colour = 16'b00000_000000_00000;
		830: oled_colour = 16'b00000_000000_00000;
		831: oled_colour = 16'b00000_000000_00000;
		832: oled_colour = 16'b00000_000000_00000;
		833: oled_colour = 16'b00000_000000_00000;
		834: oled_colour = 16'b00000_000000_00000;
		835: oled_colour = 16'b00000_000000_00000;
		836: oled_colour = 16'b00000_000000_00000;
		837: oled_colour = 16'b00000_000000_00000;
		838: oled_colour = 16'b00000_000000_00000;
		839: oled_colour = 16'b00000_000000_00000;
		840: oled_colour = 16'b00000_000000_00000;
		841: oled_colour = 16'b00000_000000_00000;
		842: oled_colour = 16'b00000_000000_00000;
		843: oled_colour = 16'b00000_000000_00000;
		844: oled_colour = 16'b00000_000000_00000;
		845: oled_colour = 16'b00000_000000_00000;
		846: oled_colour = 16'b00000_000000_00000;
		847: oled_colour = 16'b00000_000000_00000;
		848: oled_colour = 16'b00000_000000_00000;
		849: oled_colour = 16'b00000_000000_00000;
		850: oled_colour = 16'b00000_000000_00000;
		851: oled_colour = 16'b00000_000000_00000;
		852: oled_colour = 16'b00000_000000_00000;
		853: oled_colour = 16'b00000_000000_00000;
		854: oled_colour = 16'b00000_000000_00000;
		855: oled_colour = 16'b00000_000000_00000;
		856: oled_colour = 16'b00000_000000_00000;
		857: oled_colour = 16'b00000_000000_00000;
		858: oled_colour = 16'b00000_000000_00000;
		859: oled_colour = 16'b00000_000000_00000;
		860: oled_colour = 16'b00000_000000_00000;
		861: oled_colour = 16'b00000_000000_00000;
		862: oled_colour = 16'b00000_000000_00000;
		863: oled_colour = 16'b00000_000000_00000;
		864: oled_colour = 16'b00000_000000_00000;
		865: oled_colour = 16'b00000_000000_00000;
		866: oled_colour = 16'b00000_000000_00000;
		867: oled_colour = 16'b00000_000000_00000;
		868: oled_colour = 16'b00000_000000_00000;
		869: oled_colour = 16'b00000_000000_00000;
		870: oled_colour = 16'b00000_000000_00000;
		871: oled_colour = 16'b00000_000000_00000;
		872: oled_colour = 16'b00000_000000_00000;
		873: oled_colour = 16'b00000_000000_00000;
		874: oled_colour = 16'b00000_000000_00000;
		875: oled_colour = 16'b00000_000000_00000;
		876: oled_colour = 16'b00000_000000_00000;
		877: oled_colour = 16'b00000_000000_00000;
		878: oled_colour = 16'b00000_000000_00000;
		879: oled_colour = 16'b00000_000000_00000;
		880: oled_colour = 16'b00000_000000_00000;
		881: oled_colour = 16'b00000_000000_00000;
		882: oled_colour = 16'b00000_000000_00000;
		883: oled_colour = 16'b00000_000000_00000;
		884: oled_colour = 16'b00000_000000_00000;
		885: oled_colour = 16'b00000_000000_00000;
		886: oled_colour = 16'b00000_000000_00000;
		887: oled_colour = 16'b00000_000000_00000;
		888: oled_colour = 16'b00000_000000_00000;
		889: oled_colour = 16'b00000_000000_00000;
		890: oled_colour = 16'b00000_000000_00000;
		891: oled_colour = 16'b00000_000000_00000;
		892: oled_colour = 16'b00000_000000_00000;
		893: oled_colour = 16'b00000_000000_00000;
		894: oled_colour = 16'b00000_000000_00000;
		895: oled_colour = 16'b00000_000000_00000;
		896: oled_colour = 16'b00000_000000_00000;
		897: oled_colour = 16'b00000_000000_00000;
		898: oled_colour = 16'b00000_000000_00000;
		899: oled_colour = 16'b00000_000000_00000;
		900: oled_colour = 16'b00000_000000_00000;
		901: oled_colour = 16'b00000_000000_00000;
		902: oled_colour = 16'b00000_000000_00000;
		903: oled_colour = 16'b00000_000000_00000;
		904: oled_colour = 16'b00000_000000_00000;
		905: oled_colour = 16'b00000_000000_00000;
		906: oled_colour = 16'b00000_000000_00000;
		907: oled_colour = 16'b00000_000000_00000;
		908: oled_colour = 16'b00000_000000_00000;
		909: oled_colour = 16'b00000_000000_00000;
		910: oled_colour = 16'b00000_000000_00000;
		911: oled_colour = 16'b00000_000000_00000;
		912: oled_colour = 16'b00000_000000_00000;
		913: oled_colour = 16'b00000_000000_00000;
		914: oled_colour = 16'b00000_000000_00000;
		915: oled_colour = 16'b00000_000000_00000;
		916: oled_colour = 16'b00000_000000_00000;
		917: oled_colour = 16'b00000_000000_00000;
		918: oled_colour = 16'b00000_000000_00000;
		919: oled_colour = 16'b00000_000000_00000;
		920: oled_colour = 16'b00000_000000_00000;
		921: oled_colour = 16'b00000_000000_00000;
		922: oled_colour = 16'b00000_000000_00000;
		923: oled_colour = 16'b00000_000000_00000;
		924: oled_colour = 16'b00000_000000_00000;
		925: oled_colour = 16'b00000_000000_00000;
		926: oled_colour = 16'b00000_000000_00000;
		927: oled_colour = 16'b00000_000000_00000;
		928: oled_colour = 16'b00000_000000_00000;
		929: oled_colour = 16'b00000_000000_00000;
		930: oled_colour = 16'b00000_000000_00000;
		931: oled_colour = 16'b00000_000000_00000;
		932: oled_colour = 16'b00000_000000_00000;
		933: oled_colour = 16'b00000_000000_00000;
		934: oled_colour = 16'b00000_000000_00000;
		935: oled_colour = 16'b00000_000000_00000;
		936: oled_colour = 16'b00000_000000_00000;
		937: oled_colour = 16'b00000_000000_00000;
		938: oled_colour = 16'b00000_000000_00000;
		939: oled_colour = 16'b00000_000000_00000;
		940: oled_colour = 16'b00000_000000_00000;
		941: oled_colour = 16'b00000_000000_00000;
		942: oled_colour = 16'b00000_000000_00000;
		943: oled_colour = 16'b00000_000000_00000;
		944: oled_colour = 16'b00000_000000_00000;
		945: oled_colour = 16'b00000_000000_00000;
		946: oled_colour = 16'b00000_000000_00000;
		947: oled_colour = 16'b00000_000000_00000;
		948: oled_colour = 16'b00000_000000_00000;
		949: oled_colour = 16'b00000_000000_00000;
		950: oled_colour = 16'b00000_000000_00000;
		951: oled_colour = 16'b00000_000000_00000;
		952: oled_colour = 16'b00000_000000_00000;
		953: oled_colour = 16'b00000_000000_00000;
		954: oled_colour = 16'b00000_000000_00000;
		955: oled_colour = 16'b00000_000000_00000;
		956: oled_colour = 16'b00000_000000_00000;
		957: oled_colour = 16'b00000_000000_00000;
		958: oled_colour = 16'b00000_000000_00000;
		959: oled_colour = 16'b00000_000000_00000;
		960: oled_colour = 16'b00000_000000_00000;
		961: oled_colour = 16'b00000_000000_00000;
		962: oled_colour = 16'b00000_000000_00000;
		963: oled_colour = 16'b00000_000000_00000;
		964: oled_colour = 16'b00000_000000_00000;
		965: oled_colour = 16'b00000_000000_00000;
		966: oled_colour = 16'b00000_000000_00000;
		967: oled_colour = 16'b00000_000000_00000;
		968: oled_colour = 16'b00000_000000_00000;
		969: oled_colour = 16'b00000_000000_00000;
		970: oled_colour = 16'b00000_000000_00000;
		971: oled_colour = 16'b00000_000000_00000;
		972: oled_colour = 16'b00000_000000_00000;
		973: oled_colour = 16'b00000_000000_00000;
		974: oled_colour = 16'b00000_000000_00000;
		975: oled_colour = 16'b00000_000000_00000;
		976: oled_colour = 16'b00000_000000_00000;
		977: oled_colour = 16'b00000_000000_00000;
		978: oled_colour = 16'b00000_000000_00000;
		979: oled_colour = 16'b00000_000000_00000;
		980: oled_colour = 16'b00000_000000_00000;
		981: oled_colour = 16'b00000_000000_00000;
		982: oled_colour = 16'b00000_000000_00000;
		983: oled_colour = 16'b00000_000000_00000;
		984: oled_colour = 16'b00000_000000_00000;
		985: oled_colour = 16'b00000_000000_00000;
		986: oled_colour = 16'b00000_000000_00000;
		987: oled_colour = 16'b00000_000000_00000;
		988: oled_colour = 16'b00000_000000_00000;
		989: oled_colour = 16'b00000_000000_00000;
		990: oled_colour = 16'b00000_000000_00000;
		991: oled_colour = 16'b00000_000000_00000;
		992: oled_colour = 16'b00000_000000_00000;
		993: oled_colour = 16'b00000_000000_00000;
		994: oled_colour = 16'b00000_000000_00000;
		995: oled_colour = 16'b00000_000000_00000;
		996: oled_colour = 16'b00000_000000_00000;
		997: oled_colour = 16'b00000_000000_00000;
		998: oled_colour = 16'b00000_000000_00000;
		999: oled_colour = 16'b00000_000000_00000;
		1000: oled_colour = 16'b00000_000000_00000;
		1001: oled_colour = 16'b00000_000000_00000;
		1002: oled_colour = 16'b00000_000000_00000;
		1003: oled_colour = 16'b00000_000000_00000;
		1004: oled_colour = 16'b00000_000000_00000;
		1005: oled_colour = 16'b00000_000000_00000;
		1006: oled_colour = 16'b00000_000000_00000;
		1007: oled_colour = 16'b00000_000000_00000;
		1008: oled_colour = 16'b00000_000000_00000;
		1009: oled_colour = 16'b00000_000000_00000;
		1010: oled_colour = 16'b00000_000000_00000;
		1011: oled_colour = 16'b00000_000000_00000;
		1012: oled_colour = 16'b00000_000000_00000;
		1013: oled_colour = 16'b00000_000000_00000;
		1014: oled_colour = 16'b00000_000000_00000;
		1015: oled_colour = 16'b00000_000000_00000;
		1016: oled_colour = 16'b00000_000000_00000;
		1017: oled_colour = 16'b00000_000000_00000;
		1018: oled_colour = 16'b00000_000000_00000;
		1019: oled_colour = 16'b00000_000000_00000;
		1020: oled_colour = 16'b00000_000000_00000;
		1021: oled_colour = 16'b00000_000000_00000;
		1022: oled_colour = 16'b00000_000000_00000;
		1023: oled_colour = 16'b00000_000000_00000;
		1024: oled_colour = 16'b00000_000000_00000;
		1025: oled_colour = 16'b00000_000000_00000;
		1026: oled_colour = 16'b00000_000000_00000;
		1027: oled_colour = 16'b00000_000000_00000;
		1028: oled_colour = 16'b00000_000000_00000;
		1029: oled_colour = 16'b00000_000000_00000;
		1030: oled_colour = 16'b00000_000000_00000;
		1031: oled_colour = 16'b00000_000000_00000;
		1032: oled_colour = 16'b00000_000000_00000;
		1033: oled_colour = 16'b00000_000000_00000;
		1034: oled_colour = 16'b00000_000000_00000;
		1035: oled_colour = 16'b00000_000000_00000;
		1036: oled_colour = 16'b00000_000000_00000;
		1037: oled_colour = 16'b00000_000000_00000;
		1038: oled_colour = 16'b00000_000000_00000;
		1039: oled_colour = 16'b00000_000000_00000;
		1040: oled_colour = 16'b00000_000000_00000;
		1041: oled_colour = 16'b00000_000000_00000;
		1042: oled_colour = 16'b00000_000000_00000;
		1043: oled_colour = 16'b00000_000000_00000;
		1044: oled_colour = 16'b00000_000000_00000;
		1045: oled_colour = 16'b00000_000000_00000;
		1046: oled_colour = 16'b00000_000000_00000;
		1047: oled_colour = 16'b00000_000000_00000;
		1048: oled_colour = 16'b00000_000000_00000;
		1049: oled_colour = 16'b00000_000000_00000;
		1050: oled_colour = 16'b00000_000000_00000;
		1051: oled_colour = 16'b00000_000000_00000;
		1052: oled_colour = 16'b00000_000000_00000;
		1053: oled_colour = 16'b00000_000000_00000;
		1054: oled_colour = 16'b00000_000000_00000;
		1055: oled_colour = 16'b00000_000000_00000;
		1056: oled_colour = 16'b00000_000000_00000;
		1057: oled_colour = 16'b00000_000000_00000;
		1058: oled_colour = 16'b00000_000000_00000;
		1059: oled_colour = 16'b00000_000000_00000;
		1060: oled_colour = 16'b00000_000000_00000;
		1061: oled_colour = 16'b00000_000000_00000;
		1062: oled_colour = 16'b00000_000000_00000;
		1063: oled_colour = 16'b00000_000000_00000;
		1064: oled_colour = 16'b00000_000000_00000;
		1065: oled_colour = 16'b00000_000000_00000;
		1066: oled_colour = 16'b00000_000000_00000;
		1067: oled_colour = 16'b00000_000000_00000;
		1068: oled_colour = 16'b00000_000000_00000;
		1069: oled_colour = 16'b00000_000000_00000;
		1070: oled_colour = 16'b00000_000000_00000;
		1071: oled_colour = 16'b00000_000000_00000;
		1072: oled_colour = 16'b00000_000000_00000;
		1073: oled_colour = 16'b00000_000000_00000;
		1074: oled_colour = 16'b00000_000000_00000;
		1075: oled_colour = 16'b00000_000000_00000;
		1076: oled_colour = 16'b00000_000000_00000;
		1077: oled_colour = 16'b00000_000000_00000;
		1078: oled_colour = 16'b00000_000000_00000;
		1079: oled_colour = 16'b00000_000000_00000;
		1080: oled_colour = 16'b00000_000000_00000;
		1081: oled_colour = 16'b00000_000000_00000;
		1082: oled_colour = 16'b00000_000000_00000;
		1083: oled_colour = 16'b00000_000000_00000;
		1084: oled_colour = 16'b00000_000000_00000;
		1085: oled_colour = 16'b00000_000000_00000;
		1086: oled_colour = 16'b00000_000000_00000;
		1087: oled_colour = 16'b00000_000000_00000;
		1088: oled_colour = 16'b00000_000000_00000;
		1089: oled_colour = 16'b00000_000000_00000;
		1090: oled_colour = 16'b00000_000000_00000;
		1091: oled_colour = 16'b00000_000000_00000;
		1092: oled_colour = 16'b00000_000000_00000;
		1093: oled_colour = 16'b00000_000000_00000;
		1094: oled_colour = 16'b00000_000000_00000;
		1095: oled_colour = 16'b00000_000000_00000;
		1096: oled_colour = 16'b00000_000000_00000;
		1097: oled_colour = 16'b00000_000000_00000;
		1098: oled_colour = 16'b00000_000000_00000;
		1099: oled_colour = 16'b00000_000000_00000;
		1100: oled_colour = 16'b00000_000000_00000;
		1101: oled_colour = 16'b00000_000000_00000;
		1102: oled_colour = 16'b00000_000000_00000;
		1103: oled_colour = 16'b00000_000000_00000;
		1104: oled_colour = 16'b00000_000000_00000;
		1105: oled_colour = 16'b00000_000000_00000;
		1106: oled_colour = 16'b00000_000000_00000;
		1107: oled_colour = 16'b00000_000000_00000;
		1108: oled_colour = 16'b00000_000000_00000;
		1109: oled_colour = 16'b00000_000000_00000;
		1110: oled_colour = 16'b00000_000000_00000;
		1111: oled_colour = 16'b00000_000000_00000;
		1112: oled_colour = 16'b00000_000000_00000;
		1113: oled_colour = 16'b00000_000000_00000;
		1114: oled_colour = 16'b00000_000000_00000;
		1115: oled_colour = 16'b00000_000000_00000;
		1116: oled_colour = 16'b00000_000000_00000;
		1117: oled_colour = 16'b00000_000000_00000;
		1118: oled_colour = 16'b00000_000000_00000;
		1119: oled_colour = 16'b00000_000000_00000;
		1120: oled_colour = 16'b00000_000000_00000;
		1121: oled_colour = 16'b00000_000000_00000;
		1122: oled_colour = 16'b00000_000000_00000;
		1123: oled_colour = 16'b00000_000000_00000;
		1124: oled_colour = 16'b00000_000000_00000;
		1125: oled_colour = 16'b00000_000000_00000;
		1126: oled_colour = 16'b00000_000000_00000;
		1127: oled_colour = 16'b00000_000000_00000;
		1128: oled_colour = 16'b00000_000000_00000;
		1129: oled_colour = 16'b00000_000000_00000;
		1130: oled_colour = 16'b00000_000000_00000;
		1131: oled_colour = 16'b00000_000000_00000;
		1132: oled_colour = 16'b00000_000000_00000;
		1133: oled_colour = 16'b00000_000000_00000;
		1134: oled_colour = 16'b00000_000000_00000;
		1135: oled_colour = 16'b00000_000000_00000;
		1136: oled_colour = 16'b00000_000000_00000;
		1137: oled_colour = 16'b00000_000000_00000;
		1138: oled_colour = 16'b00000_000000_00000;
		1139: oled_colour = 16'b00000_000000_00000;
		1140: oled_colour = 16'b00000_000000_00000;
		1141: oled_colour = 16'b00000_000000_00000;
		1142: oled_colour = 16'b00000_000000_00000;
		1143: oled_colour = 16'b00000_000000_00000;
		1144: oled_colour = 16'b00000_000000_00000;
		1145: oled_colour = 16'b00000_000000_00000;
		1146: oled_colour = 16'b00000_000000_00000;
		1147: oled_colour = 16'b00000_000000_00000;
		1148: oled_colour = 16'b00000_000000_00000;
		1149: oled_colour = 16'b00000_000000_00000;
		1150: oled_colour = 16'b00000_000000_00000;
		1151: oled_colour = 16'b00000_000000_00000;
		1152: oled_colour = 16'b00000_000000_00000;
		1153: oled_colour = 16'b00000_000000_00000;
		1154: oled_colour = 16'b00000_000000_00000;
		1155: oled_colour = 16'b00000_000000_00000;
		1156: oled_colour = 16'b00000_000000_00000;
		1157: oled_colour = 16'b00000_000000_00000;
		1158: oled_colour = 16'b00000_000000_00000;
		1159: oled_colour = 16'b00000_000000_00000;
		1160: oled_colour = 16'b00000_000000_00000;
		1161: oled_colour = 16'b00000_000000_00000;
		1162: oled_colour = 16'b00000_000000_00000;
		1163: oled_colour = 16'b00000_000000_00000;
		1164: oled_colour = 16'b00000_000000_00000;
		1165: oled_colour = 16'b00000_000000_00000;
		1166: oled_colour = 16'b00000_000000_00000;
		1167: oled_colour = 16'b00000_000000_00000;
		1168: oled_colour = 16'b00000_000000_00000;
		1169: oled_colour = 16'b00000_000000_00000;
		1170: oled_colour = 16'b00000_000000_00000;
		1171: oled_colour = 16'b00000_000000_00000;
		1172: oled_colour = 16'b00000_000000_00000;
		1173: oled_colour = 16'b00000_000000_00000;
		1174: oled_colour = 16'b00000_000000_00000;
		1175: oled_colour = 16'b00000_000000_00000;
		1176: oled_colour = 16'b00000_000000_00000;
		1177: oled_colour = 16'b00000_000000_00000;
		1178: oled_colour = 16'b00000_000000_00000;
		1179: oled_colour = 16'b00000_000000_00000;
		1180: oled_colour = 16'b00000_000000_00000;
		1181: oled_colour = 16'b00000_000000_00000;
		1182: oled_colour = 16'b00000_000000_00000;
		1183: oled_colour = 16'b00000_000000_00000;
		1184: oled_colour = 16'b00000_000000_00000;
		1185: oled_colour = 16'b00000_000000_00000;
		1186: oled_colour = 16'b00000_000000_00000;
		1187: oled_colour = 16'b00000_000000_00000;
		1188: oled_colour = 16'b00000_000000_00000;
		1189: oled_colour = 16'b00000_000000_00000;
		1190: oled_colour = 16'b00000_000000_00000;
		1191: oled_colour = 16'b00000_000000_00000;
		1192: oled_colour = 16'b00000_000000_00000;
		1193: oled_colour = 16'b00000_000000_00000;
		1194: oled_colour = 16'b00000_000000_00000;
		1195: oled_colour = 16'b00000_000000_00000;
		1196: oled_colour = 16'b00000_000000_00000;
		1197: oled_colour = 16'b00000_000000_00000;
		1198: oled_colour = 16'b00000_000000_00000;
		1199: oled_colour = 16'b00000_000000_00000;
		1200: oled_colour = 16'b00000_000000_00000;
		1201: oled_colour = 16'b00000_000000_00000;
		1202: oled_colour = 16'b00000_000000_00000;
		1203: oled_colour = 16'b00000_000000_00000;
		1204: oled_colour = 16'b00000_000000_00000;
		1205: oled_colour = 16'b00000_000000_00000;
		1206: oled_colour = 16'b00000_000000_00000;
		1207: oled_colour = 16'b00000_000000_00000;
		1208: oled_colour = 16'b00000_000000_00000;
		1209: oled_colour = 16'b00000_000000_00000;
		1210: oled_colour = 16'b00000_000000_00000;
		1211: oled_colour = 16'b00000_000000_00000;
		1212: oled_colour = 16'b00000_000000_00000;
		1213: oled_colour = 16'b00000_000000_00000;
		1214: oled_colour = 16'b00000_000000_00000;
		1215: oled_colour = 16'b00000_000000_00000;
		1216: oled_colour = 16'b00000_000000_00000;
		1217: oled_colour = 16'b00000_000000_00000;
		1218: oled_colour = 16'b00000_000000_00000;
		1219: oled_colour = 16'b00000_000000_00000;
		1220: oled_colour = 16'b00000_000000_00000;
		1221: oled_colour = 16'b00000_000000_00000;
		1222: oled_colour = 16'b00000_000000_00000;
		1223: oled_colour = 16'b00000_000000_00000;
		1224: oled_colour = 16'b00000_000000_00000;
		1225: oled_colour = 16'b00000_000000_00000;
		1226: oled_colour = 16'b00000_000000_00000;
		1227: oled_colour = 16'b00000_000000_00000;
		1228: oled_colour = 16'b00000_000000_00000;
		1229: oled_colour = 16'b00000_000000_00000;
		1230: oled_colour = 16'b00000_000000_00000;
		1231: oled_colour = 16'b00000_000000_00000;
		1232: oled_colour = 16'b00000_000000_00000;
		1233: oled_colour = 16'b00000_000000_00000;
		1234: oled_colour = 16'b00000_000000_00000;
		1235: oled_colour = 16'b00000_000000_00000;
		1236: oled_colour = 16'b00000_000000_00000;
		1237: oled_colour = 16'b00000_000000_00000;
		1238: oled_colour = 16'b00000_000000_00000;
		1239: oled_colour = 16'b00000_000000_00000;
		1240: oled_colour = 16'b00000_000000_00000;
		1241: oled_colour = 16'b00000_000000_00000;
		1242: oled_colour = 16'b00000_000000_00000;
		1243: oled_colour = 16'b00000_000000_00000;
		1244: oled_colour = 16'b00000_000000_00000;
		1245: oled_colour = 16'b00000_000000_00000;
		1246: oled_colour = 16'b00000_000000_00000;
		1247: oled_colour = 16'b00000_000000_00000;
		1248: oled_colour = 16'b00000_000000_00000;
		1249: oled_colour = 16'b00000_000000_00000;
		1250: oled_colour = 16'b00000_000000_00000;
		1251: oled_colour = 16'b00000_000000_00000;
		1252: oled_colour = 16'b00000_000000_00000;
		1253: oled_colour = 16'b00000_000000_00000;
		1254: oled_colour = 16'b00000_000000_00000;
		1255: oled_colour = 16'b00000_000000_00000;
		1256: oled_colour = 16'b00000_000000_00000;
		1257: oled_colour = 16'b00000_000000_00000;
		1258: oled_colour = 16'b00000_000000_00000;
		1259: oled_colour = 16'b00000_000000_00000;
		1260: oled_colour = 16'b00000_000000_00000;
		1261: oled_colour = 16'b00000_000000_00000;
		1262: oled_colour = 16'b00000_000000_00000;
		1263: oled_colour = 16'b00000_000000_00000;
		1264: oled_colour = 16'b00000_000000_00000;
		1265: oled_colour = 16'b00000_000000_00000;
		1266: oled_colour = 16'b00000_000000_00000;
		1267: oled_colour = 16'b00000_000000_00000;
		1268: oled_colour = 16'b00000_000000_00000;
		1269: oled_colour = 16'b00000_000000_00000;
		1270: oled_colour = 16'b00000_000000_00000;
		1271: oled_colour = 16'b00000_000000_00000;
		1272: oled_colour = 16'b00000_000000_00000;
		1273: oled_colour = 16'b00000_000000_00000;
		1274: oled_colour = 16'b00000_000000_00000;
		1275: oled_colour = 16'b00000_000000_00000;
		1276: oled_colour = 16'b00000_000000_00000;
		1277: oled_colour = 16'b00000_000000_00000;
		1278: oled_colour = 16'b00000_000000_00000;
		1279: oled_colour = 16'b00000_000000_00000;
		1280: oled_colour = 16'b00000_000000_00000;
		1281: oled_colour = 16'b00000_000000_00000;
		1282: oled_colour = 16'b00000_000000_00000;
		1283: oled_colour = 16'b00000_000000_00000;
		1284: oled_colour = 16'b00000_000000_00000;
		1285: oled_colour = 16'b00000_000000_00000;
		1286: oled_colour = 16'b00000_000000_00000;
		1287: oled_colour = 16'b00000_000000_00000;
		1288: oled_colour = 16'b00000_000000_00000;
		1289: oled_colour = 16'b00000_000000_00000;
		1290: oled_colour = 16'b00000_000000_00000;
		1291: oled_colour = 16'b00000_000000_00000;
		1292: oled_colour = 16'b00000_000000_00000;
		1293: oled_colour = 16'b00000_000000_00000;
		1294: oled_colour = 16'b00000_000000_00000;
		1295: oled_colour = 16'b00000_000000_00000;
		1296: oled_colour = 16'b00000_000000_00000;
		1297: oled_colour = 16'b00000_000000_00000;
		1298: oled_colour = 16'b00000_000000_00000;
		1299: oled_colour = 16'b00000_000000_00000;
		1300: oled_colour = 16'b00000_000000_00000;
		1301: oled_colour = 16'b00000_000000_00000;
		1302: oled_colour = 16'b00000_000000_00000;
		1303: oled_colour = 16'b00000_000000_00000;
		1304: oled_colour = 16'b00000_000000_00000;
		1305: oled_colour = 16'b00000_000000_00000;
		1306: oled_colour = 16'b00000_000000_00000;
		1307: oled_colour = 16'b00000_000000_00000;
		1308: oled_colour = 16'b00000_000000_00000;
		1309: oled_colour = 16'b00000_000000_00000;
		1310: oled_colour = 16'b00000_000000_00000;
		1311: oled_colour = 16'b00000_000000_00000;
		1312: oled_colour = 16'b00000_000000_00000;
		1313: oled_colour = 16'b00000_000000_00000;
		1314: oled_colour = 16'b00000_000000_00000;
		1315: oled_colour = 16'b00000_000000_00000;
		1316: oled_colour = 16'b00000_000000_00000;
		1317: oled_colour = 16'b00000_000000_00000;
		1318: oled_colour = 16'b00000_000000_00000;
		1319: oled_colour = 16'b00000_000000_00000;
		1320: oled_colour = 16'b00000_000000_00000;
		1321: oled_colour = 16'b00000_000000_00000;
		1322: oled_colour = 16'b00000_000000_00000;
		1323: oled_colour = 16'b00000_000000_00000;
		1324: oled_colour = 16'b00000_000000_00000;
		1325: oled_colour = 16'b00000_000000_00000;
		1326: oled_colour = 16'b00000_000000_00000;
		1327: oled_colour = 16'b00000_000000_00000;
		1328: oled_colour = 16'b00000_000000_00000;
		1329: oled_colour = 16'b00000_000000_00000;
		1330: oled_colour = 16'b00000_000000_00000;
		1331: oled_colour = 16'b00000_000000_00000;
		1332: oled_colour = 16'b00000_000000_00000;
		1333: oled_colour = 16'b00000_000000_00000;
		1334: oled_colour = 16'b00000_000000_00000;
		1335: oled_colour = 16'b00000_000000_00000;
		1336: oled_colour = 16'b00000_000000_00000;
		1337: oled_colour = 16'b00000_000000_00000;
		1338: oled_colour = 16'b00000_000000_00000;
		1339: oled_colour = 16'b00000_000000_00000;
		1340: oled_colour = 16'b00000_000000_00000;
		1341: oled_colour = 16'b00000_000000_00000;
		1342: oled_colour = 16'b00000_000000_00000;
		1343: oled_colour = 16'b00000_000000_00000;
		1344: oled_colour = 16'b00000_000000_00000;
		1345: oled_colour = 16'b00000_000000_00000;
		1346: oled_colour = 16'b00000_000000_00000;
		1347: oled_colour = 16'b00000_000000_00000;
		1348: oled_colour = 16'b00000_000000_00000;
		1349: oled_colour = 16'b00000_000000_00000;
		1350: oled_colour = 16'b00000_000000_00000;
		1351: oled_colour = 16'b00000_000000_00000;
		1352: oled_colour = 16'b00000_000000_00000;
		1353: oled_colour = 16'b00000_000000_00000;
		1354: oled_colour = 16'b00000_000000_00000;
		1355: oled_colour = 16'b00000_000000_00000;
		1356: oled_colour = 16'b00000_000000_00000;
		1357: oled_colour = 16'b00000_000000_00000;
		1358: oled_colour = 16'b00000_000000_00000;
		1359: oled_colour = 16'b00000_000000_00000;
		1360: oled_colour = 16'b00000_000000_00000;
		1361: oled_colour = 16'b00000_000000_00000;
		1362: oled_colour = 16'b00000_000000_00000;
		1363: oled_colour = 16'b00000_000000_00000;
		1364: oled_colour = 16'b00000_000000_00000;
		1365: oled_colour = 16'b00000_000000_00000;
		1366: oled_colour = 16'b00000_000000_00000;
		1367: oled_colour = 16'b00000_000000_00000;
		1368: oled_colour = 16'b00000_000000_00000;
		1369: oled_colour = 16'b00000_000000_00000;
		1370: oled_colour = 16'b00000_000000_00000;
		1371: oled_colour = 16'b00000_000000_00000;
		1372: oled_colour = 16'b00000_000000_00000;
		1373: oled_colour = 16'b00000_000000_00000;
		1374: oled_colour = 16'b00000_000000_00000;
		1375: oled_colour = 16'b00000_000000_00000;
		1376: oled_colour = 16'b00000_000000_00000;
		1377: oled_colour = 16'b00000_000000_00000;
		1378: oled_colour = 16'b00000_000000_00000;
		1379: oled_colour = 16'b00000_000000_00000;
		1380: oled_colour = 16'b00000_000000_00000;
		1381: oled_colour = 16'b00000_000000_00000;
		1382: oled_colour = 16'b00000_000000_00000;
		1383: oled_colour = 16'b00000_000000_00000;
		1384: oled_colour = 16'b00000_000000_00000;
		1385: oled_colour = 16'b00000_000000_00000;
		1386: oled_colour = 16'b00000_000000_00000;
		1387: oled_colour = 16'b00000_000000_00000;
		1388: oled_colour = 16'b00000_000000_00000;
		1389: oled_colour = 16'b00000_000000_00000;
		1390: oled_colour = 16'b00000_000000_00000;
		1391: oled_colour = 16'b00000_000000_00000;
		1392: oled_colour = 16'b00000_000000_00000;
		1393: oled_colour = 16'b00000_000000_00000;
		1394: oled_colour = 16'b00000_000000_00000;
		1395: oled_colour = 16'b00000_000000_00000;
		1396: oled_colour = 16'b00000_000000_00000;
		1397: oled_colour = 16'b00000_000000_00000;
		1398: oled_colour = 16'b00000_000000_00000;
		1399: oled_colour = 16'b00000_000000_00000;
		1400: oled_colour = 16'b00000_000000_00000;
		1401: oled_colour = 16'b00000_000000_00000;
		1402: oled_colour = 16'b00000_000000_00000;
		1403: oled_colour = 16'b00000_000000_00000;
		1404: oled_colour = 16'b00000_000000_00000;
		1405: oled_colour = 16'b00000_000000_00000;
		1406: oled_colour = 16'b00000_000000_00000;
		1407: oled_colour = 16'b00000_000000_00000;
		1408: oled_colour = 16'b00000_000000_00000;
		1409: oled_colour = 16'b00000_000000_00000;
		1410: oled_colour = 16'b00000_000000_00000;
		1411: oled_colour = 16'b00000_000000_00000;
		1412: oled_colour = 16'b00000_000000_00000;
		1413: oled_colour = 16'b00000_000000_00000;
		1414: oled_colour = 16'b00000_000000_00000;
		1415: oled_colour = 16'b00000_000000_00000;
		1416: oled_colour = 16'b00000_000000_00000;
		1417: oled_colour = 16'b00000_000000_00000;
		1418: oled_colour = 16'b00000_000000_00000;
		1419: oled_colour = 16'b00000_000000_00000;
		1420: oled_colour = 16'b00000_000000_00000;
		1421: oled_colour = 16'b00000_000000_00000;
		1422: oled_colour = 16'b00000_000000_00000;
		1423: oled_colour = 16'b00000_000000_00000;
		1424: oled_colour = 16'b00000_000000_00000;
		1425: oled_colour = 16'b00000_000000_00000;
		1426: oled_colour = 16'b00000_000000_00000;
		1427: oled_colour = 16'b00000_000000_00000;
		1428: oled_colour = 16'b00000_000000_00000;
		1429: oled_colour = 16'b00000_000000_00000;
		1430: oled_colour = 16'b00000_000000_00000;
		1431: oled_colour = 16'b00000_000000_00000;
		1432: oled_colour = 16'b00000_000000_00000;
		1433: oled_colour = 16'b00000_000000_00000;
		1434: oled_colour = 16'b00000_000000_00000;
		1435: oled_colour = 16'b00000_000000_00000;
		1436: oled_colour = 16'b00000_000000_00000;
		1437: oled_colour = 16'b00000_000000_00000;
		1438: oled_colour = 16'b00000_000000_00000;
		1439: oled_colour = 16'b00000_000000_00000;
		1440: oled_colour = 16'b00000_000000_00000;
		1441: oled_colour = 16'b00000_000000_00000;
		1442: oled_colour = 16'b00000_000000_00000;
		1443: oled_colour = 16'b00000_000000_00000;
		1444: oled_colour = 16'b00000_000000_00000;
		1445: oled_colour = 16'b00000_000000_00000;
		1446: oled_colour = 16'b00000_000000_00000;
		1447: oled_colour = 16'b00000_000000_00000;
		1448: oled_colour = 16'b00000_000000_00000;
		1449: oled_colour = 16'b00000_000000_00000;
		1450: oled_colour = 16'b00000_000000_00000;
		1451: oled_colour = 16'b00000_000000_00000;
		1452: oled_colour = 16'b00000_000000_00000;
		1453: oled_colour = 16'b00000_000000_00000;
		1454: oled_colour = 16'b00000_000000_00000;
		1455: oled_colour = 16'b00000_000000_00000;
		1456: oled_colour = 16'b00000_000000_00000;
		1457: oled_colour = 16'b00000_000000_00000;
		1458: oled_colour = 16'b00000_000000_00000;
		1459: oled_colour = 16'b00000_000000_00000;
		1460: oled_colour = 16'b00000_000000_00000;
		1461: oled_colour = 16'b00000_000000_00000;
		1462: oled_colour = 16'b00000_000000_00000;
		1463: oled_colour = 16'b00000_000000_00000;
		1464: oled_colour = 16'b00000_000000_00000;
		1465: oled_colour = 16'b00000_000000_00000;
		1466: oled_colour = 16'b00000_000000_00000;
		1467: oled_colour = 16'b00000_000000_00000;
		1468: oled_colour = 16'b00000_000000_00000;
		1469: oled_colour = 16'b00000_000000_00000;
		1470: oled_colour = 16'b00000_000000_00000;
		1471: oled_colour = 16'b00000_000000_00000;
		1472: oled_colour = 16'b00000_000000_00000;
		1473: oled_colour = 16'b00000_000000_00000;
		1474: oled_colour = 16'b00000_000000_00000;
		1475: oled_colour = 16'b00000_000000_00000;
		1476: oled_colour = 16'b00000_000000_00000;
		1477: oled_colour = 16'b00000_000000_00000;
		1478: oled_colour = 16'b00000_000000_00000;
		1479: oled_colour = 16'b00000_000000_00000;
		1480: oled_colour = 16'b00000_000000_00000;
		1481: oled_colour = 16'b00000_000000_00000;
		1482: oled_colour = 16'b00000_000000_00000;
		1483: oled_colour = 16'b00000_000000_00000;
		1484: oled_colour = 16'b00000_000000_00000;
		1485: oled_colour = 16'b00000_000000_00000;
		1486: oled_colour = 16'b00000_000000_00000;
		1487: oled_colour = 16'b00000_000000_00000;
		1488: oled_colour = 16'b00000_000000_00000;
		1489: oled_colour = 16'b00000_000000_00000;
		1490: oled_colour = 16'b00000_000000_00000;
		1491: oled_colour = 16'b00000_000000_00000;
		1492: oled_colour = 16'b00000_000000_00000;
		1493: oled_colour = 16'b00000_000000_00000;
		1494: oled_colour = 16'b00000_000000_00000;
		1495: oled_colour = 16'b00000_000000_00000;
		1496: oled_colour = 16'b00000_000000_00000;
		1497: oled_colour = 16'b00000_000000_00000;
		1498: oled_colour = 16'b00000_000000_00000;
		1499: oled_colour = 16'b00000_000000_00000;
		1500: oled_colour = 16'b00000_000000_00000;
		1501: oled_colour = 16'b00000_000000_00000;
		1502: oled_colour = 16'b00000_000000_00000;
		1503: oled_colour = 16'b00000_000000_00000;
		1504: oled_colour = 16'b00000_000000_00000;
		1505: oled_colour = 16'b00000_000000_00000;
		1506: oled_colour = 16'b00000_000000_00000;
		1507: oled_colour = 16'b00000_000000_00000;
		1508: oled_colour = 16'b00000_000000_00000;
		1509: oled_colour = 16'b00000_000000_00000;
		1510: oled_colour = 16'b00000_000000_00000;
		1511: oled_colour = 16'b00000_000000_00000;
		1512: oled_colour = 16'b00000_000000_00000;
		1513: oled_colour = 16'b00000_000000_00000;
		1514: oled_colour = 16'b00000_000000_00000;
		1515: oled_colour = 16'b00000_000000_00000;
		1516: oled_colour = 16'b00000_000000_00000;
		1517: oled_colour = 16'b00000_000000_00000;
		1518: oled_colour = 16'b00000_000000_00000;
		1519: oled_colour = 16'b00000_000000_00000;
		1520: oled_colour = 16'b00000_000000_00000;
		1521: oled_colour = 16'b00000_000000_00000;
		1522: oled_colour = 16'b00000_000000_00000;
		1523: oled_colour = 16'b00000_000000_00000;
		1524: oled_colour = 16'b00000_000000_00000;
		1525: oled_colour = 16'b00000_000000_00000;
		1526: oled_colour = 16'b00000_000000_00000;
		1527: oled_colour = 16'b00000_000000_00000;
		1528: oled_colour = 16'b00000_000000_00000;
		1529: oled_colour = 16'b00000_000000_00000;
		1530: oled_colour = 16'b00000_000000_00000;
		1531: oled_colour = 16'b00000_000000_00000;
		1532: oled_colour = 16'b00000_000000_00000;
		1533: oled_colour = 16'b00000_000000_00000;
		1534: oled_colour = 16'b00000_000000_00000;
		1535: oled_colour = 16'b00000_000000_00000;
		1536: oled_colour = 16'b00000_000000_00000;
		1537: oled_colour = 16'b00000_000000_00000;
		1538: oled_colour = 16'b00000_000000_00000;
		1539: oled_colour = 16'b00000_000000_00000;
		1540: oled_colour = 16'b00000_000000_00000;
		1541: oled_colour = 16'b00000_000000_00000;
		1542: oled_colour = 16'b00000_000000_00000;
		1543: oled_colour = 16'b00000_000000_00000;
		1544: oled_colour = 16'b00000_000000_00000;
		1545: oled_colour = 16'b00000_000000_00000;
		1546: oled_colour = 16'b00000_000000_00000;
		1547: oled_colour = 16'b00000_000000_00000;
		1548: oled_colour = 16'b00000_000000_00000;
		1549: oled_colour = 16'b00000_000000_00000;
		1550: oled_colour = 16'b00000_000000_00000;
		1551: oled_colour = 16'b00000_000000_00000;
		1552: oled_colour = 16'b00000_000000_00000;
		1553: oled_colour = 16'b00000_000000_00000;
		1554: oled_colour = 16'b00000_000000_00000;
		1555: oled_colour = 16'b00000_000000_00000;
		1556: oled_colour = 16'b00000_000000_00000;
		1557: oled_colour = 16'b00000_000000_00000;
		1558: oled_colour = 16'b00000_000000_00000;
		1559: oled_colour = 16'b00000_000000_00000;
		1560: oled_colour = 16'b00000_000000_00000;
		1561: oled_colour = 16'b00000_000000_00000;
		1562: oled_colour = 16'b00000_000000_00000;
		1563: oled_colour = 16'b00000_000000_00000;
		1564: oled_colour = 16'b00000_000000_00000;
		1565: oled_colour = 16'b00000_000000_00000;
		1566: oled_colour = 16'b00000_000000_00000;
		1567: oled_colour = 16'b00000_000000_00000;
		1568: oled_colour = 16'b00000_000000_00000;
		1569: oled_colour = 16'b00000_000000_00000;
		1570: oled_colour = 16'b00000_000000_00000;
		1571: oled_colour = 16'b00000_000000_00000;
		1572: oled_colour = 16'b00000_000000_00000;
		1573: oled_colour = 16'b00000_000000_00000;
		1574: oled_colour = 16'b00000_000000_00000;
		1575: oled_colour = 16'b00000_000000_00000;
		1576: oled_colour = 16'b00000_000000_00000;
		1577: oled_colour = 16'b00000_000000_00000;
		1578: oled_colour = 16'b00000_000000_00000;
		1579: oled_colour = 16'b00000_000000_00000;
		1580: oled_colour = 16'b00000_000000_00000;
		1581: oled_colour = 16'b00000_000000_00000;
		1582: oled_colour = 16'b00000_000000_00000;
		1583: oled_colour = 16'b00000_000000_00000;
		1584: oled_colour = 16'b00000_000000_00000;
		1585: oled_colour = 16'b00000_000000_00000;
		1586: oled_colour = 16'b00000_000000_00000;
		1587: oled_colour = 16'b00000_000000_00000;
		1588: oled_colour = 16'b00000_000000_00000;
		1589: oled_colour = 16'b00000_000000_00000;
		1590: oled_colour = 16'b00000_000000_00000;
		1591: oled_colour = 16'b00000_000000_00000;
		1592: oled_colour = 16'b00000_000000_00000;
		1593: oled_colour = 16'b00000_000000_00000;
		1594: oled_colour = 16'b00000_000000_00000;
		1595: oled_colour = 16'b00000_000000_00000;
		1596: oled_colour = 16'b00000_000000_00000;
		1597: oled_colour = 16'b00000_000000_00000;
		1598: oled_colour = 16'b00000_000000_00000;
		1599: oled_colour = 16'b00000_000000_00000;
		1600: oled_colour = 16'b00000_000000_00000;
		1601: oled_colour = 16'b00000_000000_00000;
		1602: oled_colour = 16'b00000_000000_00000;
		1603: oled_colour = 16'b00000_000000_00000;
		1604: oled_colour = 16'b00000_000000_00000;
		1605: oled_colour = 16'b00000_000000_00000;
		1606: oled_colour = 16'b00000_000000_00000;
		1607: oled_colour = 16'b00000_000000_00000;
		1608: oled_colour = 16'b00000_000000_00000;
		1609: oled_colour = 16'b00000_000000_00000;
		1610: oled_colour = 16'b00000_000000_00000;
		1611: oled_colour = 16'b00000_000000_00000;
		1612: oled_colour = 16'b00000_000000_00000;
		1613: oled_colour = 16'b00000_000000_00000;
		1614: oled_colour = 16'b00000_000000_00000;
		1615: oled_colour = 16'b00000_000000_00000;
		1616: oled_colour = 16'b00000_000000_00000;
		1617: oled_colour = 16'b00000_000000_00000;
		1618: oled_colour = 16'b00000_000000_00000;
		1619: oled_colour = 16'b00000_000000_00000;
		1620: oled_colour = 16'b00000_000000_00000;
		1621: oled_colour = 16'b00000_000000_00000;
		1622: oled_colour = 16'b00000_000000_00000;
		1623: oled_colour = 16'b00000_000000_00000;
		1624: oled_colour = 16'b00000_000000_00000;
		1625: oled_colour = 16'b00000_000000_00000;
		1626: oled_colour = 16'b00000_000000_00000;
		1627: oled_colour = 16'b00000_000000_00000;
		1628: oled_colour = 16'b00000_000000_00000;
		1629: oled_colour = 16'b00000_000000_00000;
		1630: oled_colour = 16'b00000_000000_00000;
		1631: oled_colour = 16'b00000_000000_00000;
		1632: oled_colour = 16'b00000_000000_00000;
		1633: oled_colour = 16'b00000_000000_00000;
		1634: oled_colour = 16'b00000_000000_00000;
		1635: oled_colour = 16'b00000_000000_00000;
		1636: oled_colour = 16'b00000_000000_00000;
		1637: oled_colour = 16'b00000_000000_00000;
		1638: oled_colour = 16'b00000_000000_00000;
		1639: oled_colour = 16'b00000_000000_00000;
		1640: oled_colour = 16'b00000_000000_00000;
		1641: oled_colour = 16'b00000_000000_00000;
		1642: oled_colour = 16'b00000_000000_00000;
		1643: oled_colour = 16'b00000_000000_00000;
		1644: oled_colour = 16'b00000_000000_00000;
		1645: oled_colour = 16'b00000_000000_00000;
		1646: oled_colour = 16'b00000_000000_00000;
		1647: oled_colour = 16'b00000_000000_00000;
		1648: oled_colour = 16'b00000_000000_00000;
		1649: oled_colour = 16'b00000_000000_00000;
		1650: oled_colour = 16'b00000_000000_00000;
		1651: oled_colour = 16'b00000_000000_00000;
		1652: oled_colour = 16'b00000_000000_00000;
		1653: oled_colour = 16'b00000_000000_00000;
		1654: oled_colour = 16'b00000_000000_00000;
		1655: oled_colour = 16'b00000_000000_00000;
		1656: oled_colour = 16'b00000_000000_00000;
		1657: oled_colour = 16'b00000_000000_00000;
		1658: oled_colour = 16'b00000_000000_00000;
		1659: oled_colour = 16'b00000_000000_00000;
		1660: oled_colour = 16'b00000_000000_00000;
		1661: oled_colour = 16'b00000_000000_00000;
		1662: oled_colour = 16'b00000_000000_00000;
		1663: oled_colour = 16'b00000_000000_00000;
		1664: oled_colour = 16'b00000_000000_00000;
		1665: oled_colour = 16'b00000_000000_00000;
		1666: oled_colour = 16'b00000_000000_00000;
		1667: oled_colour = 16'b00000_000000_00000;
		1668: oled_colour = 16'b00000_000000_00000;
		1669: oled_colour = 16'b00000_000000_00000;
		1670: oled_colour = 16'b00000_000000_00000;
		1671: oled_colour = 16'b00000_000000_00000;
		1672: oled_colour = 16'b00000_000000_00000;
		1673: oled_colour = 16'b00000_000000_00000;
		1674: oled_colour = 16'b00000_000000_00000;
		1675: oled_colour = 16'b00000_000000_00000;
		1676: oled_colour = 16'b00000_000000_00000;
		1677: oled_colour = 16'b00000_000000_00000;
		1678: oled_colour = 16'b00000_000000_00000;
		1679: oled_colour = 16'b00000_000000_00000;
		1680: oled_colour = 16'b11111_111111_11111; 
		1681: oled_colour = 16'b11111_111111_11111; 
		1682: oled_colour = 16'b11111_111111_11111; 
		1683: oled_colour = 16'b11111_111111_11111; 
		1684: oled_colour = 16'b11111_111111_11111; 
		1685: oled_colour = 16'b11111_111111_11111; 
		1686: oled_colour = 16'b11111_111111_11111; 
		1687: oled_colour = 16'b11111_111111_11111; 
		1688: oled_colour = 16'b11111_111111_11111; 
		1689: oled_colour = 16'b00000_000000_00000;
		1690: oled_colour = 16'b00000_000000_00000;
		1691: oled_colour = 16'b00000_000000_00000;
		1692: oled_colour = 16'b00000_000000_00000;
		1693: oled_colour = 16'b00000_000000_00000;
		1694: oled_colour = 16'b00000_000000_00000;
		1695: oled_colour = 16'b00000_000000_00000;
		1696: oled_colour = 16'b00000_000000_00000;
		1697: oled_colour = 16'b00000_000000_00000;
		1698: oled_colour = 16'b00000_000000_00000;
		1699: oled_colour = 16'b00000_000000_00000;
		1700: oled_colour = 16'b00000_000000_00000;
		1701: oled_colour = 16'b00000_000000_00000;
		1702: oled_colour = 16'b00000_000000_00000;
		1703: oled_colour = 16'b00000_000000_00000;
		1704: oled_colour = 16'b00000_000000_00000;
		1705: oled_colour = 16'b00000_000000_00000;
		1706: oled_colour = 16'b00000_000000_00000;
		1707: oled_colour = 16'b00000_000000_00000;
		1708: oled_colour = 16'b00000_000000_00000;
		1709: oled_colour = 16'b00000_000000_00000;
		1710: oled_colour = 16'b00000_000000_00000;
		1711: oled_colour = 16'b00000_000000_00000;
		1712: oled_colour = 16'b00000_000000_00000;
		1713: oled_colour = 16'b00000_000000_00000;
		1714: oled_colour = 16'b00000_000000_00000;
		1715: oled_colour = 16'b00000_000000_00000;
		1716: oled_colour = 16'b00000_000000_00000;
		1717: oled_colour = 16'b00000_000000_00000;
		1718: oled_colour = 16'b00000_000000_00000;
		1719: oled_colour = 16'b00000_000000_00000;
		1720: oled_colour = 16'b00000_000000_00000;
		1721: oled_colour = 16'b00000_000000_00000;
		1722: oled_colour = 16'b00000_000000_00000;
		1723: oled_colour = 16'b00000_000000_00000;
		1724: oled_colour = 16'b00000_000000_00000;
		1725: oled_colour = 16'b00000_000000_00000;
		1726: oled_colour = 16'b00000_000000_00000;
		1727: oled_colour = 16'b00000_000000_00000;
		1728: oled_colour = 16'b00000_000000_00000;
		1729: oled_colour = 16'b00000_000000_00000;
		1730: oled_colour = 16'b00000_000000_00000;
		1731: oled_colour = 16'b00000_000000_00000;
		1732: oled_colour = 16'b00000_000000_00000;
		1733: oled_colour = 16'b00000_000000_00000;
		1734: oled_colour = 16'b00000_000000_00000;
		1735: oled_colour = 16'b00000_000000_00000;
		1736: oled_colour = 16'b00000_000000_00000;
		1737: oled_colour = 16'b00000_000000_00000;
		1738: oled_colour = 16'b00000_000000_00000;
		1739: oled_colour = 16'b00000_000000_00000;
		1740: oled_colour = 16'b00000_000000_00000;
		1741: oled_colour = 16'b00000_000000_00000;
		1742: oled_colour = 16'b00000_000000_00000;
		1743: oled_colour = 16'b00000_000000_00000;
		1744: oled_colour = 16'b00000_000000_00000;
		1745: oled_colour = 16'b00000_000000_00000;
		1746: oled_colour = 16'b00000_000000_00000;
		1747: oled_colour = 16'b00000_000000_00000;
		1748: oled_colour = 16'b00000_000000_00000;
		1749: oled_colour = 16'b00000_000000_00000;
		1750: oled_colour = 16'b00000_000000_00000;
		1751: oled_colour = 16'b00000_000000_00000;
		1752: oled_colour = 16'b00000_000000_00000;
		1753: oled_colour = 16'b00000_000000_00000;
		1754: oled_colour = 16'b00000_000000_00000;
		1755: oled_colour = 16'b00000_000000_00000;
		1756: oled_colour = 16'b00000_000000_00000;
		1757: oled_colour = 16'b00000_000000_00000;
		1758: oled_colour = 16'b00000_000000_00000;
		1759: oled_colour = 16'b00000_000000_00000;
		1760: oled_colour = 16'b00000_000000_00000;
		1761: oled_colour = 16'b00000_000000_00000;
		1762: oled_colour = 16'b00000_000000_00000;
		1763: oled_colour = 16'b00000_000000_00000;
		1764: oled_colour = 16'b00000_000000_00000;
		1765: oled_colour = 16'b00000_000000_00000;
		1766: oled_colour = 16'b00000_000000_00000;
		1767: oled_colour = 16'b00000_000000_00000;
		1768: oled_colour = 16'b00000_000000_00000;
		1769: oled_colour = 16'b00000_000000_00000;
		1770: oled_colour = 16'b00000_000000_00000;
		1771: oled_colour = 16'b00000_000000_00000;
		1772: oled_colour = 16'b00000_000000_00000;
		1773: oled_colour = 16'b00000_000000_00000;
		1774: oled_colour = 16'b11111_111111_11111; 
		1775: oled_colour = 16'b00000_000000_00000;
		1776: oled_colour = 16'b00000_000000_00000;
		1777: oled_colour = 16'b00000_000000_00000;
		1778: oled_colour = 16'b00000_000000_00000;
		1779: oled_colour = 16'b00000_000000_00000;
		1780: oled_colour = 16'b00000_000000_00000;
		1781: oled_colour = 16'b00000_000000_00000;
		1782: oled_colour = 16'b00000_000000_00000;
		1783: oled_colour = 16'b00000_000000_00000;
		1784: oled_colour = 16'b00000_000000_00000;
		1785: oled_colour = 16'b00000_000000_00000;
		1786: oled_colour = 16'b00000_000000_00000;
		1787: oled_colour = 16'b00000_000000_00000;
		1788: oled_colour = 16'b00000_000000_00000;
		1789: oled_colour = 16'b00000_000000_00000;
		1790: oled_colour = 16'b00000_000000_00000;
		1791: oled_colour = 16'b00000_000000_00000;
		1792: oled_colour = 16'b00000_000000_00000;
		1793: oled_colour = 16'b00000_000000_00000;
		1794: oled_colour = 16'b00000_000000_00000;
		1795: oled_colour = 16'b00000_000000_00000;
		1796: oled_colour = 16'b00000_000000_00000;
		1797: oled_colour = 16'b00000_000000_00000;
		1798: oled_colour = 16'b00000_000000_00000;
		1799: oled_colour = 16'b00000_000000_00000;
		1800: oled_colour = 16'b00000_000000_00000;
		1801: oled_colour = 16'b00000_000000_00000;
		1802: oled_colour = 16'b00000_000000_00000;
		1803: oled_colour = 16'b00000_000000_00000;
		1804: oled_colour = 16'b00000_000000_00000;
		1805: oled_colour = 16'b00000_000000_00000;
		1806: oled_colour = 16'b00000_000000_00000;
		1807: oled_colour = 16'b00000_000000_00000;
		1808: oled_colour = 16'b00000_000000_00000;
		1809: oled_colour = 16'b00000_000000_00000;
		1810: oled_colour = 16'b00000_000000_00000;
		1811: oled_colour = 16'b00000_000000_00000;
		1812: oled_colour = 16'b00000_000000_00000;
		1813: oled_colour = 16'b00000_000000_00000;
		1814: oled_colour = 16'b00000_000000_00000;
		1815: oled_colour = 16'b00000_000000_00000;
		1816: oled_colour = 16'b00000_000000_00000;
		1817: oled_colour = 16'b00000_000000_00000;
		1818: oled_colour = 16'b00000_000000_00000;
		1819: oled_colour = 16'b00000_000000_00000;
		1820: oled_colour = 16'b00000_000000_00000;
		1821: oled_colour = 16'b00000_000000_00000;
		1822: oled_colour = 16'b00000_000000_00000;
		1823: oled_colour = 16'b00000_000000_00000;
		1824: oled_colour = 16'b00000_000000_00000;
		1825: oled_colour = 16'b00000_000000_00000;
		1826: oled_colour = 16'b00000_000000_00000;
		1827: oled_colour = 16'b00000_000000_00000;
		1828: oled_colour = 16'b00000_000000_00000;
		1829: oled_colour = 16'b00000_000000_00000;
		1830: oled_colour = 16'b00000_000000_00000;
		1831: oled_colour = 16'b00000_000000_00000;
		1832: oled_colour = 16'b00000_000000_00000;
		1833: oled_colour = 16'b00000_000000_00000;
		1834: oled_colour = 16'b00000_000000_00000;
		1835: oled_colour = 16'b00000_000000_00000;
		1836: oled_colour = 16'b00000_000000_00000;
		1837: oled_colour = 16'b00000_000000_00000;
		1838: oled_colour = 16'b00000_000000_00000;
		1839: oled_colour = 16'b00000_000000_00000;
		1840: oled_colour = 16'b00000_000000_00000;
		1841: oled_colour = 16'b00000_000000_00000;
		1842: oled_colour = 16'b00000_000000_00000;
		1843: oled_colour = 16'b00000_000000_00000;
		1844: oled_colour = 16'b00000_000000_00000;
		1845: oled_colour = 16'b00000_000000_00000;
		1846: oled_colour = 16'b00000_000000_00000;
		1847: oled_colour = 16'b00000_000000_00000;
		1848: oled_colour = 16'b00000_000000_00000;
		1849: oled_colour = 16'b00000_000000_00000;
		1850: oled_colour = 16'b00000_000000_00000;
		1851: oled_colour = 16'b00000_000000_00000;
		1852: oled_colour = 16'b00000_000000_00000;
		1853: oled_colour = 16'b00000_000000_00000;
		1854: oled_colour = 16'b00000_000000_00000;
		1855: oled_colour = 16'b00000_000000_00000;
		1856: oled_colour = 16'b00000_000000_00000;
		1857: oled_colour = 16'b00000_000000_00000;
		1858: oled_colour = 16'b00000_000000_00000;
		1859: oled_colour = 16'b00000_000000_00000;
		1860: oled_colour = 16'b00000_000000_00000;
		1861: oled_colour = 16'b00000_000000_00000;
		1862: oled_colour = 16'b00000_000000_00000;
		1863: oled_colour = 16'b00000_000000_00000;
		1864: oled_colour = 16'b00000_000000_00000;
		1865: oled_colour = 16'b00000_000000_00000;
		1866: oled_colour = 16'b00000_000000_00000;
		1867: oled_colour = 16'b00000_000000_00000;
		1868: oled_colour = 16'b11111_111111_11111; 
		1869: oled_colour = 16'b00000_000000_00000;
		1870: oled_colour = 16'b00000_000000_00000;
		1871: oled_colour = 16'b11111_111111_11111; 
		1872: oled_colour = 16'b11110_111001_11100; 
		1873: oled_colour = 16'b11110_111000_11010; 
		1874: oled_colour = 16'b11111_111100_11100; 
		1875: oled_colour = 16'b11111_111101_11001; 
		1876: oled_colour = 16'b11111_111110_11001; 
		1877: oled_colour = 16'b11111_111101_11010; 
		1878: oled_colour = 16'b11111_111101_11011; 
		1879: oled_colour = 16'b11111_111110_11101; 
		1880: oled_colour = 16'b11111_111110_11101; 
		1881: oled_colour = 16'b11111_111110_11111; 
		1882: oled_colour = 16'b00000_000000_00000;
		1883: oled_colour = 16'b00000_000000_00000;
		1884: oled_colour = 16'b00000_000000_00000;
		1885: oled_colour = 16'b00000_000000_00000;
		1886: oled_colour = 16'b00000_000000_00000;
		1887: oled_colour = 16'b00000_000000_00000;
		1888: oled_colour = 16'b00000_000000_00000;
		1889: oled_colour = 16'b00000_000000_00000;
		1890: oled_colour = 16'b00000_000000_00000;
		1891: oled_colour = 16'b00000_000000_00000;
		1892: oled_colour = 16'b00000_000000_00000;
		1893: oled_colour = 16'b00000_000000_00000;
		1894: oled_colour = 16'b00000_000000_00000;
		1895: oled_colour = 16'b00000_000000_00000;
		1896: oled_colour = 16'b00000_000000_00000;
		1897: oled_colour = 16'b00000_000000_00000;
		1898: oled_colour = 16'b00000_000000_00000;
		1899: oled_colour = 16'b00000_000000_00000;
		1900: oled_colour = 16'b00000_000000_00000;
		1901: oled_colour = 16'b00000_000000_00000;
		1902: oled_colour = 16'b00000_000000_00000;
		1903: oled_colour = 16'b00000_000000_00000;
		1904: oled_colour = 16'b00000_000000_00000;
		1905: oled_colour = 16'b00000_000000_00000;
		1906: oled_colour = 16'b00000_000000_00000;
		1907: oled_colour = 16'b00000_000000_00000;
		1908: oled_colour = 16'b00000_000000_00000;
		1909: oled_colour = 16'b00000_000000_00000;
		1910: oled_colour = 16'b00000_000000_00000;
		1911: oled_colour = 16'b00000_000000_00000;
		1912: oled_colour = 16'b00000_000000_00000;
		1913: oled_colour = 16'b00000_000000_00000;
		1914: oled_colour = 16'b00000_000000_00000;
		1915: oled_colour = 16'b00000_000000_00000;
		1916: oled_colour = 16'b00000_000000_00000;
		1917: oled_colour = 16'b00000_000000_00000;
		1918: oled_colour = 16'b00000_000000_00000;
		1919: oled_colour = 16'b00000_000000_00000;
		1920: oled_colour = 16'b00000_000000_00000;
		1921: oled_colour = 16'b00000_000000_00000;
		1922: oled_colour = 16'b00000_000000_00000;
		1923: oled_colour = 16'b00000_000000_00000;
		1924: oled_colour = 16'b00000_000000_00000;
		1925: oled_colour = 16'b00000_000000_00000;
		1926: oled_colour = 16'b00000_000000_00000;
		1927: oled_colour = 16'b00000_000000_00000;
		1928: oled_colour = 16'b00000_000000_00000;
		1929: oled_colour = 16'b00000_000000_00000;
		1930: oled_colour = 16'b00000_000000_00000;
		1931: oled_colour = 16'b00000_000000_00000;
		1932: oled_colour = 16'b00000_000000_00000;
		1933: oled_colour = 16'b00000_000000_00000;
		1934: oled_colour = 16'b00000_000000_00000;
		1935: oled_colour = 16'b00000_000000_00000;
		1936: oled_colour = 16'b00000_000000_00000;
		1937: oled_colour = 16'b00000_000000_00000;
		1938: oled_colour = 16'b00000_000000_00000;
		1939: oled_colour = 16'b00000_000000_00000;
		1940: oled_colour = 16'b00000_000000_00000;
		1941: oled_colour = 16'b00000_000000_00000;
		1942: oled_colour = 16'b00000_000000_00000;
		1943: oled_colour = 16'b00000_000000_00000;
		1944: oled_colour = 16'b00000_000000_00000;
		1945: oled_colour = 16'b00000_000000_00000;
		1946: oled_colour = 16'b00000_000000_00000;
		1947: oled_colour = 16'b00000_000000_00000;
		1948: oled_colour = 16'b00000_000000_00000;
		1949: oled_colour = 16'b00000_000000_00000;
		1950: oled_colour = 16'b00000_000000_00000;
		1951: oled_colour = 16'b00000_000000_00000;
		1952: oled_colour = 16'b00000_000000_00000;
		1953: oled_colour = 16'b00000_000000_00000;
		1954: oled_colour = 16'b00000_000000_00000;
		1955: oled_colour = 16'b00000_000000_00000;
		1956: oled_colour = 16'b00000_000000_00000;
		1957: oled_colour = 16'b00000_000000_00000;
		1958: oled_colour = 16'b00000_000000_00000;
		1959: oled_colour = 16'b00000_000000_00000;
		1960: oled_colour = 16'b00000_000000_00000;
		1961: oled_colour = 16'b00000_000000_00000;
		1962: oled_colour = 16'b00000_000000_00000;
		1963: oled_colour = 16'b00000_000000_00000;
		1964: oled_colour = 16'b00000_000000_00000;
		1965: oled_colour = 16'b11111_111110_11111; 
		1966: oled_colour = 16'b11111_111101_11110; 
		1967: oled_colour = 16'b00000_000000_00000;
		1968: oled_colour = 16'b11111_111111_11111; 
		1969: oled_colour = 16'b11110_110100_10101; 
		1970: oled_colour = 16'b11101_101110_01011; 
		1971: oled_colour = 16'b11110_110101_01010; 
		1972: oled_colour = 16'b11101_110100_00101; 
		1973: oled_colour = 16'b11110_110100_01010; 
		1974: oled_colour = 16'b11110_110010_00111; 
		1975: oled_colour = 16'b11110_110100_01101; 
		1976: oled_colour = 16'b11111_111001_11000; 
		1977: oled_colour = 16'b11111_111100_11110; 
		1978: oled_colour = 16'b11111_111111_11111; 
		1979: oled_colour = 16'b00000_000000_00000;
		1980: oled_colour = 16'b00000_000000_00000;
		1981: oled_colour = 16'b00000_000000_00000;
		1982: oled_colour = 16'b00000_000000_00000;
		1983: oled_colour = 16'b00000_000000_00000;
		1984: oled_colour = 16'b00000_000000_00000;
		1985: oled_colour = 16'b00000_000000_00000;
		1986: oled_colour = 16'b00000_000000_00000;
		1987: oled_colour = 16'b00000_000000_00000;
		1988: oled_colour = 16'b00000_000000_00000;
		1989: oled_colour = 16'b00000_000000_00000;
		1990: oled_colour = 16'b00000_000000_00000;
		1991: oled_colour = 16'b00000_000000_00000;
		1992: oled_colour = 16'b00000_000000_00000;
		1993: oled_colour = 16'b00000_000000_00000;
		1994: oled_colour = 16'b00000_000000_00000;
		1995: oled_colour = 16'b00000_000000_00000;
		1996: oled_colour = 16'b00000_000000_00000;
		1997: oled_colour = 16'b00000_000000_00000;
		1998: oled_colour = 16'b00000_000000_00000;
		1999: oled_colour = 16'b00000_000000_00000;
		2000: oled_colour = 16'b00000_000000_00000;
		2001: oled_colour = 16'b00000_000000_00000;
		2002: oled_colour = 16'b00000_000000_00000;
		2003: oled_colour = 16'b00000_000000_00000;
		2004: oled_colour = 16'b00000_000000_00000;
		2005: oled_colour = 16'b00000_000000_00000;
		2006: oled_colour = 16'b00000_000000_00000;
		2007: oled_colour = 16'b00000_000000_00000;
		2008: oled_colour = 16'b00000_000000_00000;
		2009: oled_colour = 16'b00000_000000_00000;
		2010: oled_colour = 16'b00000_000000_00000;
		2011: oled_colour = 16'b00000_000000_00000;
		2012: oled_colour = 16'b00000_000000_00000;
		2013: oled_colour = 16'b00000_000000_00000;
		2014: oled_colour = 16'b00000_000000_00000;
		2015: oled_colour = 16'b00000_000000_00000;
		2016: oled_colour = 16'b00000_000000_00000;
		2017: oled_colour = 16'b00000_000000_00000;
		2018: oled_colour = 16'b00000_000000_00000;
		2019: oled_colour = 16'b00000_000000_00000;
		2020: oled_colour = 16'b00000_000000_00000;
		2021: oled_colour = 16'b00000_000000_00000;
		2022: oled_colour = 16'b00000_000000_00000;
		2023: oled_colour = 16'b00000_000000_00000;
		2024: oled_colour = 16'b00000_000000_00000;
		2025: oled_colour = 16'b00000_000000_00000;
		2026: oled_colour = 16'b00000_000000_00000;
		2027: oled_colour = 16'b00000_000000_00000;
		2028: oled_colour = 16'b00000_000000_00000;
		2029: oled_colour = 16'b00000_000000_00000;
		2030: oled_colour = 16'b00000_000000_00000;
		2031: oled_colour = 16'b00000_000000_00000;
		2032: oled_colour = 16'b00000_000000_00000;
		2033: oled_colour = 16'b00000_000000_00000;
		2034: oled_colour = 16'b00000_000000_00000;
		2035: oled_colour = 16'b00000_000000_00000;
		2036: oled_colour = 16'b00000_000000_00000;
		2037: oled_colour = 16'b00000_000000_00000;
		2038: oled_colour = 16'b00000_000000_00000;
		2039: oled_colour = 16'b00000_000000_00000;
		2040: oled_colour = 16'b00000_000000_00000;
		2041: oled_colour = 16'b00000_000000_00000;
		2042: oled_colour = 16'b00000_000000_00000;
		2043: oled_colour = 16'b00000_000000_00000;
		2044: oled_colour = 16'b00000_000000_00000;
		2045: oled_colour = 16'b00000_000000_00000;
		2046: oled_colour = 16'b00000_000000_00000;
		2047: oled_colour = 16'b00000_000000_00000;
		2048: oled_colour = 16'b00000_000000_00000;
		2049: oled_colour = 16'b00000_000000_00000;
		2050: oled_colour = 16'b00000_000000_00000;
		2051: oled_colour = 16'b00000_000000_00000;
		2052: oled_colour = 16'b00000_000000_00000;
		2053: oled_colour = 16'b00000_000000_00000;
		2054: oled_colour = 16'b00000_000000_00000;
		2055: oled_colour = 16'b00000_000000_00000;
		2056: oled_colour = 16'b00000_000000_00000;
		2057: oled_colour = 16'b00000_000000_00000;
		2058: oled_colour = 16'b11111_111111_11111; 
		2059: oled_colour = 16'b11111_111111_11111; 
		2060: oled_colour = 16'b11101_110101_11010; 
		2061: oled_colour = 16'b11011_101101_10011; 
		2062: oled_colour = 16'b11101_110011_11000; 
		2063: oled_colour = 16'b11011_110001_10101; 
		2064: oled_colour = 16'b10111_110000_10101; 
		2065: oled_colour = 16'b11001_101011_10100; 
		2066: oled_colour = 16'b11010_100111_01100; 
		2067: oled_colour = 16'b11101_110000_01100; 
		2068: oled_colour = 16'b11100_101111_10010; 
		2069: oled_colour = 16'b11101_110001_01111; 
		2070: oled_colour = 16'b11101_110010_10011; 
		2071: oled_colour = 16'b11111_111111_11111; 
		2072: oled_colour = 16'b00000_000000_00000;
		2073: oled_colour = 16'b00000_000000_00000;
		2074: oled_colour = 16'b00000_000000_00000;
		2075: oled_colour = 16'b11111_111111_11111; 
		2076: oled_colour = 16'b00000_000000_00000;
		2077: oled_colour = 16'b00000_000000_00000;
		2078: oled_colour = 16'b00000_000000_00000;
		2079: oled_colour = 16'b00000_000000_00000;
		2080: oled_colour = 16'b00000_000000_00000;
		2081: oled_colour = 16'b00000_000000_00000;
		2082: oled_colour = 16'b00000_000000_00000;
		2083: oled_colour = 16'b00000_000000_00000;
		2084: oled_colour = 16'b00000_000000_00000;
		2085: oled_colour = 16'b00000_000000_00000;
		2086: oled_colour = 16'b00000_000000_00000;
		2087: oled_colour = 16'b00000_000000_00000;
		2088: oled_colour = 16'b00000_000000_00000;
		2089: oled_colour = 16'b00000_000000_00000;
		2090: oled_colour = 16'b00000_000000_00000;
		2091: oled_colour = 16'b00000_000000_00000;
		2092: oled_colour = 16'b00000_000000_00000;
		2093: oled_colour = 16'b00000_000000_00000;
		2094: oled_colour = 16'b00000_000000_00000;
		2095: oled_colour = 16'b00000_000000_00000;
		2096: oled_colour = 16'b00000_000000_00000;
		2097: oled_colour = 16'b00000_000000_00000;
		2098: oled_colour = 16'b00000_000000_00000;
		2099: oled_colour = 16'b00000_000000_00000;
		2100: oled_colour = 16'b00000_000000_00000;
		2101: oled_colour = 16'b00000_000000_00000;
		2102: oled_colour = 16'b00000_000000_00000;
		2103: oled_colour = 16'b00000_000000_00000;
		2104: oled_colour = 16'b00000_000000_00000;
		2105: oled_colour = 16'b00000_000000_00000;
		2106: oled_colour = 16'b00000_000000_00000;
		2107: oled_colour = 16'b00000_000000_00000;
		2108: oled_colour = 16'b00000_000000_00000;
		2109: oled_colour = 16'b00000_000000_00000;
		2110: oled_colour = 16'b00000_000000_00000;
		2111: oled_colour = 16'b00000_000000_00000;
		2112: oled_colour = 16'b00000_000000_00000;
		2113: oled_colour = 16'b00000_000000_00000;
		2114: oled_colour = 16'b00000_000000_00000;
		2115: oled_colour = 16'b00000_000000_00000;
		2116: oled_colour = 16'b00000_000000_00000;
		2117: oled_colour = 16'b00000_000000_00000;
		2118: oled_colour = 16'b00000_000000_00000;
		2119: oled_colour = 16'b00000_000000_00000;
		2120: oled_colour = 16'b00000_000000_00000;
		2121: oled_colour = 16'b00000_000000_00000;
		2122: oled_colour = 16'b00000_000000_00000;
		2123: oled_colour = 16'b00000_000000_00000;
		2124: oled_colour = 16'b00000_000000_00000;
		2125: oled_colour = 16'b00000_000000_00000;
		2126: oled_colour = 16'b00000_000000_00000;
		2127: oled_colour = 16'b00000_000000_00000;
		2128: oled_colour = 16'b00000_000000_00000;
		2129: oled_colour = 16'b00000_000000_00000;
		2130: oled_colour = 16'b00000_000000_00000;
		2131: oled_colour = 16'b00000_000000_00000;
		2132: oled_colour = 16'b00000_000000_00000;
		2133: oled_colour = 16'b00000_000000_00000;
		2134: oled_colour = 16'b00000_000000_00000;
		2135: oled_colour = 16'b00000_000000_00000;
		2136: oled_colour = 16'b00000_000000_00000;
		2137: oled_colour = 16'b00000_000000_00000;
		2138: oled_colour = 16'b00000_000000_00000;
		2139: oled_colour = 16'b00000_000000_00000;
		2140: oled_colour = 16'b00000_000000_00000;
		2141: oled_colour = 16'b00000_000000_00000;
		2142: oled_colour = 16'b00000_000000_00000;
		2143: oled_colour = 16'b00000_000000_00000;
		2144: oled_colour = 16'b00000_000000_00000;
		2145: oled_colour = 16'b00000_000000_00000;
		2146: oled_colour = 16'b00000_000000_00000;
		2147: oled_colour = 16'b00000_000000_00000;
		2148: oled_colour = 16'b00000_000000_00000;
		2149: oled_colour = 16'b00000_000000_00000;
		2150: oled_colour = 16'b00000_000000_00000;
		2151: oled_colour = 16'b00000_000000_00000;
		2152: oled_colour = 16'b00000_000000_00000;
		2153: oled_colour = 16'b11111_111111_11111; 
		2154: oled_colour = 16'b00000_000000_00000;
		2155: oled_colour = 16'b11111_111101_11110; 
		2156: oled_colour = 16'b11010_101010_10010; 
		2157: oled_colour = 16'b11101_101111_10011; 
		2158: oled_colour = 16'b11101_110011_10110; 
		2159: oled_colour = 16'b11100_101011_10000; 
		2160: oled_colour = 16'b01110_100001_01001; 
		2161: oled_colour = 16'b01110_010111_00101; 
		2162: oled_colour = 16'b11001_100110_10000; 
		2163: oled_colour = 16'b11010_100111_01110; 
		2164: oled_colour = 16'b11011_101100_10100; 
		2165: oled_colour = 16'b11001_101001_10011; 
		2166: oled_colour = 16'b11011_101100_10011; 
		2167: oled_colour = 16'b11111_111110_11111; 
		2168: oled_colour = 16'b11111_111100_11110; 
		2169: oled_colour = 16'b11011_110000_10111; 
		2170: oled_colour = 16'b11110_111001_11100; 
		2171: oled_colour = 16'b00000_000000_00000;
		2172: oled_colour = 16'b11111_111111_11111; 
		2173: oled_colour = 16'b00000_000000_00000;
		2174: oled_colour = 16'b00000_000000_00000;
		2175: oled_colour = 16'b00000_000000_00000;
		2176: oled_colour = 16'b00000_000000_00000;
		2177: oled_colour = 16'b00000_000000_00000;
		2178: oled_colour = 16'b00000_000000_00000;
		2179: oled_colour = 16'b00000_000000_00000;
		2180: oled_colour = 16'b00000_000000_00000;
		2181: oled_colour = 16'b00000_000000_00000;
		2182: oled_colour = 16'b00000_000000_00000;
		2183: oled_colour = 16'b00000_000000_00000;
		2184: oled_colour = 16'b00000_000000_00000;
		2185: oled_colour = 16'b00000_000000_00000;
		2186: oled_colour = 16'b00000_000000_00000;
		2187: oled_colour = 16'b00000_000000_00000;
		2188: oled_colour = 16'b00000_000000_00000;
		2189: oled_colour = 16'b00000_000000_00000;
		2190: oled_colour = 16'b00000_000000_00000;
		2191: oled_colour = 16'b00000_000000_00000;
		2192: oled_colour = 16'b00000_000000_00000;
		2193: oled_colour = 16'b00000_000000_00000;
		2194: oled_colour = 16'b00000_000000_00000;
		2195: oled_colour = 16'b00000_000000_00000;
		2196: oled_colour = 16'b00000_000000_00000;
		2197: oled_colour = 16'b00000_000000_00000;
		2198: oled_colour = 16'b00000_000000_00000;
		2199: oled_colour = 16'b00000_000000_00000;
		2200: oled_colour = 16'b00000_000000_00000;
		2201: oled_colour = 16'b00000_000000_00000;
		2202: oled_colour = 16'b00000_000000_00000;
		2203: oled_colour = 16'b00000_000000_00000;
		2204: oled_colour = 16'b00000_000000_00000;
		2205: oled_colour = 16'b00000_000000_00000;
		2206: oled_colour = 16'b00000_000000_00000;
		2207: oled_colour = 16'b00000_000000_00000;
		2208: oled_colour = 16'b00000_000000_00000;
		2209: oled_colour = 16'b00000_000000_00000;
		2210: oled_colour = 16'b00000_000000_00000;
		2211: oled_colour = 16'b00000_000000_00000;
		2212: oled_colour = 16'b00000_000000_00000;
		2213: oled_colour = 16'b00000_000000_00000;
		2214: oled_colour = 16'b00000_000000_00000;
		2215: oled_colour = 16'b00000_000000_00000;
		2216: oled_colour = 16'b00000_000000_00000;
		2217: oled_colour = 16'b00000_000000_00000;
		2218: oled_colour = 16'b00000_000000_00000;
		2219: oled_colour = 16'b00000_000000_00000;
		2220: oled_colour = 16'b00000_000000_00000;
		2221: oled_colour = 16'b00000_000000_00000;
		2222: oled_colour = 16'b00000_000000_00000;
		2223: oled_colour = 16'b00000_000000_00000;
		2224: oled_colour = 16'b00000_000000_00000;
		2225: oled_colour = 16'b00000_000000_00000;
		2226: oled_colour = 16'b00000_000000_00000;
		2227: oled_colour = 16'b00000_000000_00000;
		2228: oled_colour = 16'b00000_000000_00000;
		2229: oled_colour = 16'b00000_000000_00000;
		2230: oled_colour = 16'b00000_000000_00000;
		2231: oled_colour = 16'b00000_000000_00000;
		2232: oled_colour = 16'b00000_000000_00000;
		2233: oled_colour = 16'b00000_000000_00000;
		2234: oled_colour = 16'b00000_000000_00000;
		2235: oled_colour = 16'b00000_000000_00000;
		2236: oled_colour = 16'b00000_000000_00000;
		2237: oled_colour = 16'b00000_000000_00000;
		2238: oled_colour = 16'b00000_000000_00000;
		2239: oled_colour = 16'b00000_000000_00000;
		2240: oled_colour = 16'b00000_000000_00000;
		2241: oled_colour = 16'b00000_000000_00000;
		2242: oled_colour = 16'b00000_000000_00000;
		2243: oled_colour = 16'b00000_000000_00000;
		2244: oled_colour = 16'b00000_000000_00000;
		2245: oled_colour = 16'b00000_000000_00000;
		2246: oled_colour = 16'b00000_000000_00000;
		2247: oled_colour = 16'b00000_000000_00000;
		2248: oled_colour = 16'b00000_000000_00000;
		2249: oled_colour = 16'b11111_111111_11111; 
		2250: oled_colour = 16'b00000_000000_00000;
		2251: oled_colour = 16'b11101_111011_11101; 
		2252: oled_colour = 16'b10110_100001_01100; 
		2253: oled_colour = 16'b10111_011101_01011; 
		2254: oled_colour = 16'b10111_100100_10001; 
		2255: oled_colour = 16'b11011_101001_10001; 
		2256: oled_colour = 16'b10011_011101_01011; 
		2257: oled_colour = 16'b10110_011111_01011; 
		2258: oled_colour = 16'b11111_101101_10011; 
		2259: oled_colour = 16'b11001_100110_01111; 
		2260: oled_colour = 16'b11011_101100_10011; 
		2261: oled_colour = 16'b11000_101010_10001; 
		2262: oled_colour = 16'b11011_101100_10001; 
		2263: oled_colour = 16'b11110_110101_11010; 
		2264: oled_colour = 16'b11010_101111_10110; 
		2265: oled_colour = 16'b10110_100001_01100; 
		2266: oled_colour = 16'b10111_100010_01110; 
		2267: oled_colour = 16'b11110_110111_11011; 
		2268: oled_colour = 16'b00000_000000_00000;
		2269: oled_colour = 16'b11111_111111_11111; 
		2270: oled_colour = 16'b00000_000000_00000;
		2271: oled_colour = 16'b00000_000000_00000;
		2272: oled_colour = 16'b00000_000000_00000;
		2273: oled_colour = 16'b00000_000000_00000;
		2274: oled_colour = 16'b00000_000000_00000;
		2275: oled_colour = 16'b00000_000000_00000;
		2276: oled_colour = 16'b00000_000000_00000;
		2277: oled_colour = 16'b00000_000000_00000;
		2278: oled_colour = 16'b00000_000000_00000;
		2279: oled_colour = 16'b00000_000000_00000;
		2280: oled_colour = 16'b00000_000000_00000;
		2281: oled_colour = 16'b00000_000000_00000;
		2282: oled_colour = 16'b00000_000000_00000;
		2283: oled_colour = 16'b00000_000000_00000;
		2284: oled_colour = 16'b00000_000000_00000;
		2285: oled_colour = 16'b00000_000000_00000;
		2286: oled_colour = 16'b00000_000000_00000;
		2287: oled_colour = 16'b00000_000000_00000;
		2288: oled_colour = 16'b00000_000000_00000;
		2289: oled_colour = 16'b00000_000000_00000;
		2290: oled_colour = 16'b00000_000000_00000;
		2291: oled_colour = 16'b00000_000000_00000;
		2292: oled_colour = 16'b00000_000000_00000;
		2293: oled_colour = 16'b00000_000000_00000;
		2294: oled_colour = 16'b00000_000000_00000;
		2295: oled_colour = 16'b00000_000000_00000;
		2296: oled_colour = 16'b00000_000000_00000;
		2297: oled_colour = 16'b00000_000000_00000;
		2298: oled_colour = 16'b00000_000000_00000;
		2299: oled_colour = 16'b00000_000000_00000;
		2300: oled_colour = 16'b00000_000000_00000;
		2301: oled_colour = 16'b00000_000000_00000;
		2302: oled_colour = 16'b00000_000000_00000;
		2303: oled_colour = 16'b00000_000000_00000;
		2304: oled_colour = 16'b00000_000000_00000;
		2305: oled_colour = 16'b00000_000000_00000;
		2306: oled_colour = 16'b00000_000000_00000;
		2307: oled_colour = 16'b00000_000000_00000;
		2308: oled_colour = 16'b00000_000000_00000;
		2309: oled_colour = 16'b00000_000000_00000;
		2310: oled_colour = 16'b00000_000000_00000;
		2311: oled_colour = 16'b00000_000000_00000;
		2312: oled_colour = 16'b00000_000000_00000;
		2313: oled_colour = 16'b00000_000000_00000;
		2314: oled_colour = 16'b00000_000000_00000;
		2315: oled_colour = 16'b00000_000000_00000;
		2316: oled_colour = 16'b00000_000000_00000;
		2317: oled_colour = 16'b00000_000000_00000;
		2318: oled_colour = 16'b00000_000000_00000;
		2319: oled_colour = 16'b00000_000000_00000;
		2320: oled_colour = 16'b00000_000000_00000;
		2321: oled_colour = 16'b00000_000000_00000;
		2322: oled_colour = 16'b00000_000000_00000;
		2323: oled_colour = 16'b00000_000000_00000;
		2324: oled_colour = 16'b00000_000000_00000;
		2325: oled_colour = 16'b00000_000000_00000;
		2326: oled_colour = 16'b00000_000000_00000;
		2327: oled_colour = 16'b00000_000000_00000;
		2328: oled_colour = 16'b00000_000000_00000;
		2329: oled_colour = 16'b00000_000000_00000;
		2330: oled_colour = 16'b00000_000000_00000;
		2331: oled_colour = 16'b00000_000000_00000;
		2332: oled_colour = 16'b00000_000000_00000;
		2333: oled_colour = 16'b00000_000000_00000;
		2334: oled_colour = 16'b00000_000000_00000;
		2335: oled_colour = 16'b00000_000000_00000;
		2336: oled_colour = 16'b00000_000000_00000;
		2337: oled_colour = 16'b00000_000000_00000;
		2338: oled_colour = 16'b00000_000000_00000;
		2339: oled_colour = 16'b00000_000000_00000;
		2340: oled_colour = 16'b00000_000000_00000;
		2341: oled_colour = 16'b00000_000000_00000;
		2342: oled_colour = 16'b00000_000000_00000;
		2343: oled_colour = 16'b00000_000000_00000;
		2344: oled_colour = 16'b00000_000000_00000;
		2345: oled_colour = 16'b11111_111111_11111; 
		2346: oled_colour = 16'b00000_000000_00000;
		2347: oled_colour = 16'b11011_111010_11100; 
		2348: oled_colour = 16'b01111_011100_00111; 
		2349: oled_colour = 16'b11101_100111_01111; 
		2350: oled_colour = 16'b11100_101100_10010; 
		2351: oled_colour = 16'b11001_101000_10000; 
		2352: oled_colour = 16'b11000_100100_01101; 
		2353: oled_colour = 16'b11110_101110_10010; 
		2354: oled_colour = 16'b11001_100110_01111; 
		2355: oled_colour = 16'b10100_011101_01010; 
		2356: oled_colour = 16'b10101_100000_01100; 
		2357: oled_colour = 16'b10011_100000_01011; 
		2358: oled_colour = 16'b11011_101100_10011; 
		2359: oled_colour = 16'b11001_101000_10001; 
		2360: oled_colour = 16'b11000_100011_01110; 
		2361: oled_colour = 16'b11001_100111_01111; 
		2362: oled_colour = 16'b10111_100010_01101; 
		2363: oled_colour = 16'b11100_110101_11010; 
		2364: oled_colour = 16'b00000_000000_00000;
		2365: oled_colour = 16'b11111_111111_11111; 
		2366: oled_colour = 16'b00000_000000_00000;
		2367: oled_colour = 16'b00000_000000_00000;
		2368: oled_colour = 16'b00000_000000_00000;
		2369: oled_colour = 16'b00000_000000_00000;
		2370: oled_colour = 16'b00000_000000_00000;
		2371: oled_colour = 16'b00000_000000_00000;
		2372: oled_colour = 16'b00000_000000_00000;
		2373: oled_colour = 16'b00000_000000_00000;
		2374: oled_colour = 16'b00000_000000_00000;
		2375: oled_colour = 16'b00000_000000_00000;
		2376: oled_colour = 16'b00000_000000_00000;
		2377: oled_colour = 16'b00000_000000_00000;
		2378: oled_colour = 16'b00000_000000_00000;
		2379: oled_colour = 16'b00000_000000_00000;
		2380: oled_colour = 16'b00000_000000_00000;
		2381: oled_colour = 16'b00000_000000_00000;
		2382: oled_colour = 16'b00000_000000_00000;
		2383: oled_colour = 16'b00000_000000_00000;
		2384: oled_colour = 16'b00000_000000_00000;
		2385: oled_colour = 16'b00000_000000_00000;
		2386: oled_colour = 16'b00000_000000_00000;
		2387: oled_colour = 16'b00000_000000_00000;
		2388: oled_colour = 16'b00000_000000_00000;
		2389: oled_colour = 16'b00000_000000_00000;
		2390: oled_colour = 16'b00000_000000_00000;
		2391: oled_colour = 16'b00000_000000_00000;
		2392: oled_colour = 16'b00000_000000_00000;
		2393: oled_colour = 16'b00000_000000_00000;
		2394: oled_colour = 16'b00000_000000_00000;
		2395: oled_colour = 16'b00000_000000_00000;
		2396: oled_colour = 16'b00000_000000_00000;
		2397: oled_colour = 16'b00000_000000_00000;
		2398: oled_colour = 16'b00000_000000_00000;
		2399: oled_colour = 16'b00000_000000_00000;
		2400: oled_colour = 16'b00000_000000_00000;
		2401: oled_colour = 16'b00000_000000_00000;
		2402: oled_colour = 16'b00000_000000_00000;
		2403: oled_colour = 16'b00000_000000_00000;
		2404: oled_colour = 16'b00000_000000_00000;
		2405: oled_colour = 16'b00000_000000_00000;
		2406: oled_colour = 16'b00000_000000_00000;
		2407: oled_colour = 16'b00000_000000_00000;
		2408: oled_colour = 16'b00000_000000_00000;
		2409: oled_colour = 16'b00000_000000_00000;
		2410: oled_colour = 16'b00000_000000_00000;
		2411: oled_colour = 16'b00000_000000_00000;
		2412: oled_colour = 16'b00000_000000_00000;
		2413: oled_colour = 16'b00000_000000_00000;
		2414: oled_colour = 16'b00000_000000_00000;
		2415: oled_colour = 16'b00000_000000_00000;
		2416: oled_colour = 16'b00000_000000_00000;
		2417: oled_colour = 16'b00000_000000_00000;
		2418: oled_colour = 16'b00000_000000_00000;
		2419: oled_colour = 16'b00000_000000_00000;
		2420: oled_colour = 16'b00000_000000_00000;
		2421: oled_colour = 16'b00000_000000_00000;
		2422: oled_colour = 16'b00000_000000_00000;
		2423: oled_colour = 16'b00000_000000_00000;
		2424: oled_colour = 16'b00000_000000_00000;
		2425: oled_colour = 16'b00000_000000_00000;
		2426: oled_colour = 16'b00000_000000_00000;
		2427: oled_colour = 16'b00000_000000_00000;
		2428: oled_colour = 16'b00000_000000_00000;
		2429: oled_colour = 16'b00000_000000_00000;
		2430: oled_colour = 16'b00000_000000_00000;
		2431: oled_colour = 16'b00000_000000_00000;
		2432: oled_colour = 16'b00000_000000_00000;
		2433: oled_colour = 16'b00000_000000_00000;
		2434: oled_colour = 16'b00000_000000_00000;
		2435: oled_colour = 16'b00000_000000_00000;
		2436: oled_colour = 16'b00000_000000_00000;
		2437: oled_colour = 16'b00000_000000_00000;
		2438: oled_colour = 16'b00000_000000_00000;
		2439: oled_colour = 16'b00000_000000_00000;
		2440: oled_colour = 16'b00000_000000_00000;
		2441: oled_colour = 16'b11111_111111_11111; 
		2442: oled_colour = 16'b00000_000000_00000;
		2443: oled_colour = 16'b11111_111110_11111; 
		2444: oled_colour = 16'b01101_011101_01001; 
		2445: oled_colour = 16'b11000_100001_01101; 
		2446: oled_colour = 16'b11001_100111_01111; 
		2447: oled_colour = 16'b11101_110101_10111; 
		2448: oled_colour = 16'b11111_111001_11000; 
		2449: oled_colour = 16'b11000_100110_01101; 
		2450: oled_colour = 16'b01100_011011_01000; 
		2451: oled_colour = 16'b10000_011110_01001; 
		2452: oled_colour = 16'b01101_011111_01001; 
		2453: oled_colour = 16'b01001_011001_00110; 
		2454: oled_colour = 16'b11001_100111_10001; 
		2455: oled_colour = 16'b11011_100110_01111; 
		2456: oled_colour = 16'b11100_101010_10000; 
		2457: oled_colour = 16'b11001_101001_10010; 
		2458: oled_colour = 16'b11111_111100_11110; 
		2459: oled_colour = 16'b00000_000000_00000;
		2460: oled_colour = 16'b00000_000000_00000;
		2461: oled_colour = 16'b00000_000000_00000;
		2462: oled_colour = 16'b00000_000000_00000;
		2463: oled_colour = 16'b00000_000000_00000;
		2464: oled_colour = 16'b00000_000000_00000;
		2465: oled_colour = 16'b00000_000000_00000;
		2466: oled_colour = 16'b00000_000000_00000;
		2467: oled_colour = 16'b00000_000000_00000;
		2468: oled_colour = 16'b00000_000000_00000;
		2469: oled_colour = 16'b00000_000000_00000;
		2470: oled_colour = 16'b00000_000000_00000;
		2471: oled_colour = 16'b00000_000000_00000;
		2472: oled_colour = 16'b00000_000000_00000;
		2473: oled_colour = 16'b00000_000000_00000;
		2474: oled_colour = 16'b00000_000000_00000;
		2475: oled_colour = 16'b00000_000000_00000;
		2476: oled_colour = 16'b00000_000000_00000;
		2477: oled_colour = 16'b00000_000000_00000;
		2478: oled_colour = 16'b00000_000000_00000;
		2479: oled_colour = 16'b00000_000000_00000;
		2480: oled_colour = 16'b00000_000000_00000;
		2481: oled_colour = 16'b00000_000000_00000;
		2482: oled_colour = 16'b00000_000000_00000;
		2483: oled_colour = 16'b00000_000000_00000;
		2484: oled_colour = 16'b00000_000000_00000;
		2485: oled_colour = 16'b00000_000000_00000;
		2486: oled_colour = 16'b00000_000000_00000;
		2487: oled_colour = 16'b00000_000000_00000;
		2488: oled_colour = 16'b00000_000000_00000;
		2489: oled_colour = 16'b00000_000000_00000;
		2490: oled_colour = 16'b00000_000000_00000;
		2491: oled_colour = 16'b00000_000000_00000;
		2492: oled_colour = 16'b00000_000000_00000;
		2493: oled_colour = 16'b00000_000000_00000;
		2494: oled_colour = 16'b00000_000000_00000;
		2495: oled_colour = 16'b00000_000000_00000;
		2496: oled_colour = 16'b00000_000000_00000;
		2497: oled_colour = 16'b00000_000000_00000;
		2498: oled_colour = 16'b00000_000000_00000;
		2499: oled_colour = 16'b00000_000000_00000;
		2500: oled_colour = 16'b00000_000000_00000;
		2501: oled_colour = 16'b00000_000000_00000;
		2502: oled_colour = 16'b00000_000000_00000;
		2503: oled_colour = 16'b00000_000000_00000;
		2504: oled_colour = 16'b00000_000000_00000;
		2505: oled_colour = 16'b00000_000000_00000;
		2506: oled_colour = 16'b00000_000000_00000;
		2507: oled_colour = 16'b00000_000000_00000;
		2508: oled_colour = 16'b00000_000000_00000;
		2509: oled_colour = 16'b00000_000000_00000;
		2510: oled_colour = 16'b00000_000000_00000;
		2511: oled_colour = 16'b00000_000000_00000;
		2512: oled_colour = 16'b00000_000000_00000;
		2513: oled_colour = 16'b00000_000000_00000;
		2514: oled_colour = 16'b00000_000000_00000;
		2515: oled_colour = 16'b00000_000000_00000;
		2516: oled_colour = 16'b00000_000000_00000;
		2517: oled_colour = 16'b00000_000000_00000;
		2518: oled_colour = 16'b00000_000000_00000;
		2519: oled_colour = 16'b00000_000000_00000;
		2520: oled_colour = 16'b00000_000000_00000;
		2521: oled_colour = 16'b00000_000000_00000;
		2522: oled_colour = 16'b00000_000000_00000;
		2523: oled_colour = 16'b00000_000000_00000;
		2524: oled_colour = 16'b00000_000000_00000;
		2525: oled_colour = 16'b00000_000000_00000;
		2526: oled_colour = 16'b00000_000000_00000;
		2527: oled_colour = 16'b00000_000000_00000;
		2528: oled_colour = 16'b00000_000000_00000;
		2529: oled_colour = 16'b00000_000000_00000;
		2530: oled_colour = 16'b00000_000000_00000;
		2531: oled_colour = 16'b00000_000000_00000;
		2532: oled_colour = 16'b00000_000000_00000;
		2533: oled_colour = 16'b00000_000000_00000;
		2534: oled_colour = 16'b00000_000000_00000;
		2535: oled_colour = 16'b00000_000000_00000;
		2536: oled_colour = 16'b00000_000000_00000;
		2537: oled_colour = 16'b00000_000000_00000;
		2538: oled_colour = 16'b11111_111111_11111; 
		2539: oled_colour = 16'b00000_000000_00000;
		2540: oled_colour = 16'b01110_100100_01101; 
		2541: oled_colour = 16'b10011_011011_01000; 
		2542: oled_colour = 16'b11111_110101_10111; 
		2543: oled_colour = 16'b11101_101111_10101; 
		2544: oled_colour = 16'b10111_011111_01011; 
		2545: oled_colour = 16'b01001_011000_00101; 
		2546: oled_colour = 16'b01000_011110_01000; 
		2547: oled_colour = 16'b00111_011011_00110; 
		2548: oled_colour = 16'b01110_100100_01101; 
		2549: oled_colour = 16'b10000_011000_00111; 
		2550: oled_colour = 16'b11010_100100_01110; 
		2551: oled_colour = 16'b11111_110110_10111; 
		2552: oled_colour = 16'b11011_101011_10001; 
		2553: oled_colour = 16'b11111_111100_11110; 
		2554: oled_colour = 16'b00000_000000_00000;
		2555: oled_colour = 16'b11111_111111_11111; 
		2556: oled_colour = 16'b00000_000000_00000;
		2557: oled_colour = 16'b00000_000000_00000;
		2558: oled_colour = 16'b00000_000000_00000;
		2559: oled_colour = 16'b00000_000000_00000;
		2560: oled_colour = 16'b00000_000000_00000;
		2561: oled_colour = 16'b00000_000000_00000;
		2562: oled_colour = 16'b00000_000000_00000;
		2563: oled_colour = 16'b00000_000000_00000;
		2564: oled_colour = 16'b00000_000000_00000;
		2565: oled_colour = 16'b00000_000000_00000;
		2566: oled_colour = 16'b00000_000000_00000;
		2567: oled_colour = 16'b00000_000000_00000;
		2568: oled_colour = 16'b00000_000000_00000;
		2569: oled_colour = 16'b00000_000000_00000;
		2570: oled_colour = 16'b00000_000000_00000;
		2571: oled_colour = 16'b00000_000000_00000;
		2572: oled_colour = 16'b00000_000000_00000;
		2573: oled_colour = 16'b00000_000000_00000;
		2574: oled_colour = 16'b00000_000000_00000;
		2575: oled_colour = 16'b00000_000000_00000;
		2576: oled_colour = 16'b00000_000000_00000;
		2577: oled_colour = 16'b00000_000000_00000;
		2578: oled_colour = 16'b00000_000000_00000;
		2579: oled_colour = 16'b00000_000000_00000;
		2580: oled_colour = 16'b00000_000000_00000;
		2581: oled_colour = 16'b00000_000000_00000;
		2582: oled_colour = 16'b00000_000000_00000;
		2583: oled_colour = 16'b00000_000000_00000;
		2584: oled_colour = 16'b00000_000000_00000;
		2585: oled_colour = 16'b00000_000000_00000;
		2586: oled_colour = 16'b00000_000000_00000;
		2587: oled_colour = 16'b00000_000000_00000;
		2588: oled_colour = 16'b00000_000000_00000;
		2589: oled_colour = 16'b00000_000000_00000;
		2590: oled_colour = 16'b00000_000000_00000;
		2591: oled_colour = 16'b00000_000000_00000;
		2592: oled_colour = 16'b00000_000000_00000;
		2593: oled_colour = 16'b00000_000000_00000;
		2594: oled_colour = 16'b00000_000000_00000;
		2595: oled_colour = 16'b00000_000000_00000;
		2596: oled_colour = 16'b00000_000000_00000;
		2597: oled_colour = 16'b00000_000000_00000;
		2598: oled_colour = 16'b00000_000000_00000;
		2599: oled_colour = 16'b00000_000000_00000;
		2600: oled_colour = 16'b00000_000000_00000;
		2601: oled_colour = 16'b00000_000000_00000;
		2602: oled_colour = 16'b00000_000000_00000;
		2603: oled_colour = 16'b00000_000000_00000;
		2604: oled_colour = 16'b00000_000000_00000;
		2605: oled_colour = 16'b00000_000000_00000;
		2606: oled_colour = 16'b00000_000000_00000;
		2607: oled_colour = 16'b00000_000000_00000;
		2608: oled_colour = 16'b00000_000000_00000;
		2609: oled_colour = 16'b00000_000000_00000;
		2610: oled_colour = 16'b00000_000000_00000;
		2611: oled_colour = 16'b00000_000000_00000;
		2612: oled_colour = 16'b00000_000000_00000;
		2613: oled_colour = 16'b00000_000000_00000;
		2614: oled_colour = 16'b00000_000000_00000;
		2615: oled_colour = 16'b00000_000000_00000;
		2616: oled_colour = 16'b00000_000000_00000;
		2617: oled_colour = 16'b00000_000000_00000;
		2618: oled_colour = 16'b00000_000000_00000;
		2619: oled_colour = 16'b00000_000000_00000;
		2620: oled_colour = 16'b00000_000000_00000;
		2621: oled_colour = 16'b00000_000000_00000;
		2622: oled_colour = 16'b00000_000000_00000;
		2623: oled_colour = 16'b00000_000000_00000;
		2624: oled_colour = 16'b00000_000000_00000;
		2625: oled_colour = 16'b00000_000000_00000;
		2626: oled_colour = 16'b00000_000000_00000;
		2627: oled_colour = 16'b00000_000000_00000;
		2628: oled_colour = 16'b00000_000000_00000;
		2629: oled_colour = 16'b00000_000000_00000;
		2630: oled_colour = 16'b00000_000000_00000;
		2631: oled_colour = 16'b00000_000000_00000;
		2632: oled_colour = 16'b00000_000000_00000;
		2633: oled_colour = 16'b00000_000000_00000;
		2634: oled_colour = 16'b11111_111111_11111; 
		2635: oled_colour = 16'b11111_111111_11111; 
		2636: oled_colour = 16'b10011_101010_10001; 
		2637: oled_colour = 16'b01110_011010_00111; 
		2638: oled_colour = 16'b11000_100110_01110; 
		2639: oled_colour = 16'b01010_010101_00011; 
		2640: oled_colour = 16'b00100_010100_00001; 
		2641: oled_colour = 16'b00001_010011_00001; 
		2642: oled_colour = 16'b00001_010011_00001; 
		2643: oled_colour = 16'b10100_101101_10011; 
		2644: oled_colour = 16'b11111_111111_11111; 
		2645: oled_colour = 16'b11011_101101_10101; 
		2646: oled_colour = 16'b11011_101100_10011; 
		2647: oled_colour = 16'b11010_101001_10001; 
		2648: oled_colour = 16'b11100_110100_11001; 
		2649: oled_colour = 16'b00000_000000_00000;
		2650: oled_colour = 16'b11111_111111_11111; 
		2651: oled_colour = 16'b00000_000000_00000;
		2652: oled_colour = 16'b00000_000000_00000;
		2653: oled_colour = 16'b00000_000000_00000;
		2654: oled_colour = 16'b00000_000000_00000;
		2655: oled_colour = 16'b00000_000000_00000;
		2656: oled_colour = 16'b00000_000000_00000;
		2657: oled_colour = 16'b00000_000000_00000;
		2658: oled_colour = 16'b00000_000000_00000;
		2659: oled_colour = 16'b00000_000000_00000;
		2660: oled_colour = 16'b00000_000000_00000;
		2661: oled_colour = 16'b00000_000000_00000;
		2662: oled_colour = 16'b00000_000000_00000;
		2663: oled_colour = 16'b00000_000000_00000;
		2664: oled_colour = 16'b00000_000000_00000;
		2665: oled_colour = 16'b00000_000000_00000;
		2666: oled_colour = 16'b00000_000000_00000;
		2667: oled_colour = 16'b00000_000000_00000;
		2668: oled_colour = 16'b00000_000000_00000;
		2669: oled_colour = 16'b00000_000000_00000;
		2670: oled_colour = 16'b00000_000000_00000;
		2671: oled_colour = 16'b00000_000000_00000;
		2672: oled_colour = 16'b00000_000000_00000;
		2673: oled_colour = 16'b00000_000000_00000;
		2674: oled_colour = 16'b00000_000000_00000;
		2675: oled_colour = 16'b00000_000000_00000;
		2676: oled_colour = 16'b00000_000000_00000;
		2677: oled_colour = 16'b00000_000000_00000;
		2678: oled_colour = 16'b00000_000000_00000;
		2679: oled_colour = 16'b00000_000000_00000;
		2680: oled_colour = 16'b00000_000000_00000;
		2681: oled_colour = 16'b00000_000000_00000;
		2682: oled_colour = 16'b00000_000000_00000;
		2683: oled_colour = 16'b00000_000000_00000;
		2684: oled_colour = 16'b00000_000000_00000;
		2685: oled_colour = 16'b00000_000000_00000;
		2686: oled_colour = 16'b00000_000000_00000;
		2687: oled_colour = 16'b00000_000000_00000;
		2688: oled_colour = 16'b00000_000000_00000;
		2689: oled_colour = 16'b00000_000000_00000;
		2690: oled_colour = 16'b00000_000000_00000;
		2691: oled_colour = 16'b00000_000000_00000;
		2692: oled_colour = 16'b00000_000000_00000;
		2693: oled_colour = 16'b00000_000000_00000;
		2694: oled_colour = 16'b00000_000000_00000;
		2695: oled_colour = 16'b00000_000000_00000;
		2696: oled_colour = 16'b00000_000000_00000;
		2697: oled_colour = 16'b00000_000000_00000;
		2698: oled_colour = 16'b00000_000000_00000;
		2699: oled_colour = 16'b00000_000000_00000;
		2700: oled_colour = 16'b00000_000000_00000;
		2701: oled_colour = 16'b00000_000000_00000;
		2702: oled_colour = 16'b00000_000000_00000;
		2703: oled_colour = 16'b00000_000000_00000;
		2704: oled_colour = 16'b00000_000000_00000;
		2705: oled_colour = 16'b00000_000000_00000;
		2706: oled_colour = 16'b00000_000000_00000;
		2707: oled_colour = 16'b00000_000000_00000;
		2708: oled_colour = 16'b00000_000000_00000;
		2709: oled_colour = 16'b00000_000000_00000;
		2710: oled_colour = 16'b00000_000000_00000;
		2711: oled_colour = 16'b00000_000000_00000;
		2712: oled_colour = 16'b00000_000000_00000;
		2713: oled_colour = 16'b00000_000000_00000;
		2714: oled_colour = 16'b00000_000000_00000;
		2715: oled_colour = 16'b00000_000000_00000;
		2716: oled_colour = 16'b00000_000000_00000;
		2717: oled_colour = 16'b00000_000000_00000;
		2718: oled_colour = 16'b00000_000000_00000;
		2719: oled_colour = 16'b00000_000000_00000;
		2720: oled_colour = 16'b00000_000000_00000;
		2721: oled_colour = 16'b00000_000000_00000;
		2722: oled_colour = 16'b00000_000000_00000;
		2723: oled_colour = 16'b00000_000000_00000;
		2724: oled_colour = 16'b00000_000000_00000;
		2725: oled_colour = 16'b00000_000000_00000;
		2726: oled_colour = 16'b00000_000000_00000;
		2727: oled_colour = 16'b00000_000000_00000;
		2728: oled_colour = 16'b00000_000000_00000;
		2729: oled_colour = 16'b00000_000000_00000;
		2730: oled_colour = 16'b11111_111111_11111; 
		2731: oled_colour = 16'b00000_000000_00000;
		2732: oled_colour = 16'b10011_100111_10000; 
		2733: oled_colour = 16'b01100_010111_00110; 
		2734: oled_colour = 16'b01110_011000_00110; 
		2735: oled_colour = 16'b01011_011010_00101; 
		2736: oled_colour = 16'b01011_011010_00101; 
		2737: oled_colour = 16'b01100_100000_01001; 
		2738: oled_colour = 16'b01010_010110_00100; 
		2739: oled_colour = 16'b11101_111000_11100; 
		2740: oled_colour = 16'b00000_000000_00000;
		2741: oled_colour = 16'b11111_111111_11111; 
		2742: oled_colour = 16'b11111_111011_11101; 
		2743: oled_colour = 16'b11111_111100_11110; 
		2744: oled_colour = 16'b00000_000000_00000;
		2745: oled_colour = 16'b11111_111111_11111; 
		2746: oled_colour = 16'b00000_000000_00000;
		2747: oled_colour = 16'b00000_000000_00000;
		2748: oled_colour = 16'b00000_000000_00000;
		2749: oled_colour = 16'b00000_000000_00000;
		2750: oled_colour = 16'b00000_000000_00000;
		2751: oled_colour = 16'b00000_000000_00000;
		2752: oled_colour = 16'b00000_000000_00000;
		2753: oled_colour = 16'b00000_000000_00000;
		2754: oled_colour = 16'b00000_000000_00000;
		2755: oled_colour = 16'b00000_000000_00000;
		2756: oled_colour = 16'b00000_000000_00000;
		2757: oled_colour = 16'b00000_000000_00000;
		2758: oled_colour = 16'b00000_000000_00000;
		2759: oled_colour = 16'b00000_000000_00000;
		2760: oled_colour = 16'b00000_000000_00000;
		2761: oled_colour = 16'b00000_000000_00000;
		2762: oled_colour = 16'b00000_000000_00000;
		2763: oled_colour = 16'b00000_000000_00000;
		2764: oled_colour = 16'b00000_000000_00000;
		2765: oled_colour = 16'b00000_000000_00000;
		2766: oled_colour = 16'b00000_000000_00000;
		2767: oled_colour = 16'b00000_000000_00000;
		2768: oled_colour = 16'b00000_000000_00000;
		2769: oled_colour = 16'b00000_000000_00000;
		2770: oled_colour = 16'b00000_000000_00000;
		2771: oled_colour = 16'b00000_000000_00000;
		2772: oled_colour = 16'b00000_000000_00000;
		2773: oled_colour = 16'b00000_000000_00000;
		2774: oled_colour = 16'b00000_000000_00000;
		2775: oled_colour = 16'b00000_000000_00000;
		2776: oled_colour = 16'b00000_000000_00000;
		2777: oled_colour = 16'b00000_000000_00000;
		2778: oled_colour = 16'b00000_000000_00000;
		2779: oled_colour = 16'b00000_000000_00000;
		2780: oled_colour = 16'b00000_000000_00000;
		2781: oled_colour = 16'b00000_000000_00000;
		2782: oled_colour = 16'b00000_000000_00000;
		2783: oled_colour = 16'b00000_000000_00000;
		2784: oled_colour = 16'b00000_000000_00000;
		2785: oled_colour = 16'b00000_000000_00000;
		2786: oled_colour = 16'b00000_000000_00000;
		2787: oled_colour = 16'b00000_000000_00000;
		2788: oled_colour = 16'b00000_000000_00000;
		2789: oled_colour = 16'b00000_000000_00000;
		2790: oled_colour = 16'b00000_000000_00000;
		2791: oled_colour = 16'b00000_000000_00000;
		2792: oled_colour = 16'b00000_000000_00000;
		2793: oled_colour = 16'b00000_000000_00000;
		2794: oled_colour = 16'b00000_000000_00000;
		2795: oled_colour = 16'b00000_000000_00000;
		2796: oled_colour = 16'b00000_000000_00000;
		2797: oled_colour = 16'b00000_000000_00000;
		2798: oled_colour = 16'b00000_000000_00000;
		2799: oled_colour = 16'b00000_000000_00000;
		2800: oled_colour = 16'b00000_000000_00000;
		2801: oled_colour = 16'b00000_000000_00000;
		2802: oled_colour = 16'b00000_000000_00000;
		2803: oled_colour = 16'b00000_000000_00000;
		2804: oled_colour = 16'b00000_000000_00000;
		2805: oled_colour = 16'b00000_000000_00000;
		2806: oled_colour = 16'b00000_000000_00000;
		2807: oled_colour = 16'b00000_000000_00000;
		2808: oled_colour = 16'b00000_000000_00000;
		2809: oled_colour = 16'b00000_000000_00000;
		2810: oled_colour = 16'b00000_000000_00000;
		2811: oled_colour = 16'b00000_000000_00000;
		2812: oled_colour = 16'b00000_000000_00000;
		2813: oled_colour = 16'b00000_000000_00000;
		2814: oled_colour = 16'b00000_000000_00000;
		2815: oled_colour = 16'b00000_000000_00000;
		2816: oled_colour = 16'b00000_000000_00000;
		2817: oled_colour = 16'b00000_000000_00000;
		2818: oled_colour = 16'b00000_000000_00000;
		2819: oled_colour = 16'b00000_000000_00000;
		2820: oled_colour = 16'b00000_000000_00000;
		2821: oled_colour = 16'b00000_000000_00000;
		2822: oled_colour = 16'b00000_000000_00000;
		2823: oled_colour = 16'b00000_000000_00000;
		2824: oled_colour = 16'b00000_000000_00000;
		2825: oled_colour = 16'b11111_111111_11111; 
		2826: oled_colour = 16'b00000_000000_00000;
		2827: oled_colour = 16'b11101_111001_11101; 
		2828: oled_colour = 16'b10011_011011_01001; 
		2829: oled_colour = 16'b10001_100100_01101; 
		2830: oled_colour = 16'b10001_011001_01000; 
		2831: oled_colour = 16'b10011_011000_01000; 
		2832: oled_colour = 16'b01110_011111_01010; 
		2833: oled_colour = 16'b01010_011101_01000; 
		2834: oled_colour = 16'b01111_010110_00101; 
		2835: oled_colour = 16'b11101_110111_11010; 
		2836: oled_colour = 16'b11111_111111_11111; 
		2837: oled_colour = 16'b11111_111111_11111; 
		2838: oled_colour = 16'b00000_000000_00000;
		2839: oled_colour = 16'b00000_000000_00000;
		2840: oled_colour = 16'b11111_111111_11111; 
		2841: oled_colour = 16'b00000_000000_00000;
		2842: oled_colour = 16'b00000_000000_00000;
		2843: oled_colour = 16'b00000_000000_00000;
		2844: oled_colour = 16'b00000_000000_00000;
		2845: oled_colour = 16'b00000_000000_00000;
		2846: oled_colour = 16'b00000_000000_00000;
		2847: oled_colour = 16'b00000_000000_00000;
		2848: oled_colour = 16'b00000_000000_00000;
		2849: oled_colour = 16'b00000_000000_00000;
		2850: oled_colour = 16'b00000_000000_00000;
		2851: oled_colour = 16'b00000_000000_00000;
		2852: oled_colour = 16'b00000_000000_00000;
		2853: oled_colour = 16'b00000_000000_00000;
		2854: oled_colour = 16'b00000_000000_00000;
		2855: oled_colour = 16'b00000_000000_00000;
		2856: oled_colour = 16'b00000_000000_00000;
		2857: oled_colour = 16'b00000_000000_00000;
		2858: oled_colour = 16'b00000_000000_00000;
		2859: oled_colour = 16'b00000_000000_00000;
		2860: oled_colour = 16'b00000_000000_00000;
		2861: oled_colour = 16'b00000_000000_00000;
		2862: oled_colour = 16'b00000_000000_00000;
		2863: oled_colour = 16'b00000_000000_00000;
		2864: oled_colour = 16'b00000_000000_00000;
		2865: oled_colour = 16'b00000_000000_00000;
		2866: oled_colour = 16'b00000_000000_00000;
		2867: oled_colour = 16'b00000_000000_00000;
		2868: oled_colour = 16'b00000_000000_00000;
		2869: oled_colour = 16'b00000_000000_00000;
		2870: oled_colour = 16'b00000_000000_00000;
		2871: oled_colour = 16'b00000_000000_00000;
		2872: oled_colour = 16'b00000_000000_00000;
		2873: oled_colour = 16'b00000_000000_00000;
		2874: oled_colour = 16'b00000_000000_00000;
		2875: oled_colour = 16'b00000_000000_00000;
		2876: oled_colour = 16'b00000_000000_00000;
		2877: oled_colour = 16'b00000_000000_00000;
		2878: oled_colour = 16'b00000_000000_00000;
		2879: oled_colour = 16'b00000_000000_00000;
		2880: oled_colour = 16'b00000_000000_00000;
		2881: oled_colour = 16'b00000_000000_00000;
		2882: oled_colour = 16'b00000_000000_00000;
		2883: oled_colour = 16'b00000_000000_00000;
		2884: oled_colour = 16'b00000_000000_00000;
		2885: oled_colour = 16'b00000_000000_00000;
		2886: oled_colour = 16'b00000_000000_00000;
		2887: oled_colour = 16'b00000_000000_00000;
		2888: oled_colour = 16'b00000_000000_00000;
		2889: oled_colour = 16'b00000_000000_00000;
		2890: oled_colour = 16'b00000_000000_00000;
		2891: oled_colour = 16'b00000_000000_00000;
		2892: oled_colour = 16'b00000_000000_00000;
		2893: oled_colour = 16'b00000_000000_00000;
		2894: oled_colour = 16'b00000_000000_00000;
		2895: oled_colour = 16'b00000_000000_00000;
		2896: oled_colour = 16'b00000_000000_00000;
		2897: oled_colour = 16'b00000_000000_00000;
		2898: oled_colour = 16'b00000_000000_00000;
		2899: oled_colour = 16'b00000_000000_00000;
		2900: oled_colour = 16'b00000_000000_00000;
		2901: oled_colour = 16'b00000_000000_00000;
		2902: oled_colour = 16'b00000_000000_00000;
		2903: oled_colour = 16'b00000_000000_00000;
		2904: oled_colour = 16'b00000_000000_00000;
		2905: oled_colour = 16'b00000_000000_00000;
		2906: oled_colour = 16'b00000_000000_00000;
		2907: oled_colour = 16'b00000_000000_00000;
		2908: oled_colour = 16'b00000_000000_00000;
		2909: oled_colour = 16'b00000_000000_00000;
		2910: oled_colour = 16'b00000_000000_00000;
		2911: oled_colour = 16'b00000_000000_00000;
		2912: oled_colour = 16'b00000_000000_00000;
		2913: oled_colour = 16'b00000_000000_00000;
		2914: oled_colour = 16'b00000_000000_00000;
		2915: oled_colour = 16'b00000_000000_00000;
		2916: oled_colour = 16'b00000_000000_00000;
		2917: oled_colour = 16'b00000_000000_00000;
		2918: oled_colour = 16'b00000_000000_00000;
		2919: oled_colour = 16'b00000_000000_00000;
		2920: oled_colour = 16'b00000_000000_00000;
		2921: oled_colour = 16'b11111_111111_11111; 
		2922: oled_colour = 16'b00000_000000_00000;
		2923: oled_colour = 16'b11011_110100_11000; 
		2924: oled_colour = 16'b10010_100100_01110; 
		2925: oled_colour = 16'b10111_110000_10010; 
		2926: oled_colour = 16'b10110_101010_10000; 
		2927: oled_colour = 16'b10001_011001_01000; 
		2928: oled_colour = 16'b01001_011000_00101; 
		2929: oled_colour = 16'b00101_011000_00100; 
		2930: oled_colour = 16'b01010_010100_00011; 
		2931: oled_colour = 16'b10111_110001_10110; 
		2932: oled_colour = 16'b00000_000000_00000;
		2933: oled_colour = 16'b11111_111111_11111; 
		2934: oled_colour = 16'b11111_111111_11111; 
		2935: oled_colour = 16'b11111_111111_11111; 
		2936: oled_colour = 16'b00000_000000_00000;
		2937: oled_colour = 16'b00000_000000_00000;
		2938: oled_colour = 16'b00000_000000_00000;
		2939: oled_colour = 16'b00000_000000_00000;
		2940: oled_colour = 16'b00000_000000_00000;
		2941: oled_colour = 16'b00000_000000_00000;
		2942: oled_colour = 16'b00000_000000_00000;
		2943: oled_colour = 16'b00000_000000_00000;
		2944: oled_colour = 16'b00000_000000_00000;
		2945: oled_colour = 16'b00000_000000_00000;
		2946: oled_colour = 16'b00000_000000_00000;
		2947: oled_colour = 16'b00000_000000_00000;
		2948: oled_colour = 16'b00000_000000_00000;
		2949: oled_colour = 16'b00000_000000_00000;
		2950: oled_colour = 16'b00000_000000_00000;
		2951: oled_colour = 16'b00000_000000_00000;
		2952: oled_colour = 16'b00000_000000_00000;
		2953: oled_colour = 16'b00000_000000_00000;
		2954: oled_colour = 16'b00000_000000_00000;
		2955: oled_colour = 16'b00000_000000_00000;
		2956: oled_colour = 16'b00000_000000_00000;
		2957: oled_colour = 16'b00000_000000_00000;
		2958: oled_colour = 16'b00000_000000_00000;
		2959: oled_colour = 16'b00000_000000_00000;
		2960: oled_colour = 16'b00000_000000_00000;
		2961: oled_colour = 16'b00000_000000_00000;
		2962: oled_colour = 16'b00000_000000_00000;
		2963: oled_colour = 16'b00000_000000_00000;
		2964: oled_colour = 16'b00000_000000_00000;
		2965: oled_colour = 16'b00000_000000_00000;
		2966: oled_colour = 16'b00000_000000_00000;
		2967: oled_colour = 16'b00000_000000_00000;
		2968: oled_colour = 16'b00000_000000_00000;
		2969: oled_colour = 16'b00000_000000_00000;
		2970: oled_colour = 16'b00000_000000_00000;
		2971: oled_colour = 16'b00000_000000_00000;
		2972: oled_colour = 16'b00000_000000_00000;
		2973: oled_colour = 16'b00000_000000_00000;
		2974: oled_colour = 16'b00000_000000_00000;
		2975: oled_colour = 16'b00000_000000_00000;
		2976: oled_colour = 16'b00000_000000_00000;
		2977: oled_colour = 16'b00000_000000_00000;
		2978: oled_colour = 16'b00000_000000_00000;
		2979: oled_colour = 16'b00000_000000_00000;
		2980: oled_colour = 16'b00000_000000_00000;
		2981: oled_colour = 16'b00000_000000_00000;
		2982: oled_colour = 16'b00000_000000_00000;
		2983: oled_colour = 16'b00000_000000_00000;
		2984: oled_colour = 16'b00000_000000_00000;
		2985: oled_colour = 16'b00000_000000_00000;
		2986: oled_colour = 16'b00000_000000_00000;
		2987: oled_colour = 16'b00000_000000_00000;
		2988: oled_colour = 16'b00000_000000_00000;
		2989: oled_colour = 16'b00000_000000_00000;
		2990: oled_colour = 16'b00000_000000_00000;
		2991: oled_colour = 16'b00000_000000_00000;
		2992: oled_colour = 16'b00000_000000_00000;
		2993: oled_colour = 16'b00000_000000_00000;
		2994: oled_colour = 16'b00000_000000_00000;
		2995: oled_colour = 16'b00000_000000_00000;
		2996: oled_colour = 16'b00000_000000_00000;
		2997: oled_colour = 16'b00000_000000_00000;
		2998: oled_colour = 16'b00000_000000_00000;
		2999: oled_colour = 16'b00000_000000_00000;
		3000: oled_colour = 16'b00000_000000_00000;
		3001: oled_colour = 16'b00000_000000_00000;
		3002: oled_colour = 16'b00000_000000_00000;
		3003: oled_colour = 16'b00000_000000_00000;
		3004: oled_colour = 16'b00000_000000_00000;
		3005: oled_colour = 16'b00000_000000_00000;
		3006: oled_colour = 16'b00000_000000_00000;
		3007: oled_colour = 16'b00000_000000_00000;
		3008: oled_colour = 16'b00000_000000_00000;
		3009: oled_colour = 16'b00000_000000_00000;
		3010: oled_colour = 16'b00000_000000_00000;
		3011: oled_colour = 16'b00000_000000_00000;
		3012: oled_colour = 16'b00000_000000_00000;
		3013: oled_colour = 16'b00000_000000_00000;
		3014: oled_colour = 16'b00000_000000_00000;
		3015: oled_colour = 16'b00000_000000_00000;
		3016: oled_colour = 16'b00000_000000_00000;
		3017: oled_colour = 16'b11111_111111_11111; 
		3018: oled_colour = 16'b00000_000000_00000;
		3019: oled_colour = 16'b11101_111100_11100; 
		3020: oled_colour = 16'b10011_101111_10011; 
		3021: oled_colour = 16'b10011_110011_10010; 
		3022: oled_colour = 16'b11010_111101_10100; 
		3023: oled_colour = 16'b10001_101100_01111; 
		3024: oled_colour = 16'b01000_011000_00100; 
		3025: oled_colour = 16'b00110_011001_00100; 
		3026: oled_colour = 16'b01010_011001_00110; 
		3027: oled_colour = 16'b10101_110000_10110; 
		3028: oled_colour = 16'b00000_000000_00000;
		3029: oled_colour = 16'b11111_111111_11111; 
		3030: oled_colour = 16'b00000_000000_00000;
		3031: oled_colour = 16'b00000_000000_00000;
		3032: oled_colour = 16'b00000_000000_00000;
		3033: oled_colour = 16'b00000_000000_00000;
		3034: oled_colour = 16'b00000_000000_00000;
		3035: oled_colour = 16'b00000_000000_00000;
		3036: oled_colour = 16'b00000_000000_00000;
		3037: oled_colour = 16'b00000_000000_00000;
		3038: oled_colour = 16'b00000_000000_00000;
		3039: oled_colour = 16'b00000_000000_00000;
		3040: oled_colour = 16'b00000_000000_00000;
		3041: oled_colour = 16'b00000_000000_00000;
		3042: oled_colour = 16'b00000_000000_00000;
		3043: oled_colour = 16'b00000_000000_00000;
		3044: oled_colour = 16'b00000_000000_00000;
		3045: oled_colour = 16'b00000_000000_00000;
		3046: oled_colour = 16'b00000_000000_00000;
		3047: oled_colour = 16'b00000_000000_00000;
		3048: oled_colour = 16'b00000_000000_00000;
		3049: oled_colour = 16'b00000_000000_00000;
		3050: oled_colour = 16'b00000_000000_00000;
		3051: oled_colour = 16'b00000_000000_00000;
		3052: oled_colour = 16'b00000_000000_00000;
		3053: oled_colour = 16'b00000_000000_00000;
		3054: oled_colour = 16'b00000_000000_00000;
		3055: oled_colour = 16'b00000_000000_00000;
		3056: oled_colour = 16'b00000_000000_00000;
		3057: oled_colour = 16'b00000_000000_00000;
		3058: oled_colour = 16'b00000_000000_00000;
		3059: oled_colour = 16'b00000_000000_00000;
		3060: oled_colour = 16'b00000_000000_00000;
		3061: oled_colour = 16'b00000_000000_00000;
		3062: oled_colour = 16'b00000_000000_00000;
		3063: oled_colour = 16'b00000_000000_00000;
		3064: oled_colour = 16'b00000_000000_00000;
		3065: oled_colour = 16'b00000_000000_00000;
		3066: oled_colour = 16'b00000_000000_00000;
		3067: oled_colour = 16'b00000_000000_00000;
		3068: oled_colour = 16'b00000_000000_00000;
		3069: oled_colour = 16'b00000_000000_00000;
		3070: oled_colour = 16'b00000_000000_00000;
		3071: oled_colour = 16'b00000_000000_00000;
		3072: oled_colour = 16'b00000_000000_00000;
		3073: oled_colour = 16'b00000_000000_00000;
		3074: oled_colour = 16'b00000_000000_00000;
		3075: oled_colour = 16'b00000_000000_00000;
		3076: oled_colour = 16'b00000_000000_00000;
		3077: oled_colour = 16'b00000_000000_00000;
		3078: oled_colour = 16'b00000_000000_00000;
		3079: oled_colour = 16'b00000_000000_00000;
		3080: oled_colour = 16'b00000_000000_00000;
		3081: oled_colour = 16'b00000_000000_00000;
		3082: oled_colour = 16'b00000_000000_00000;
		3083: oled_colour = 16'b00000_000000_00000;
		3084: oled_colour = 16'b00000_000000_00000;
		3085: oled_colour = 16'b00000_000000_00000;
		3086: oled_colour = 16'b00000_000000_00000;
		3087: oled_colour = 16'b00000_000000_00000;
		3088: oled_colour = 16'b00000_000000_00000;
		3089: oled_colour = 16'b00000_000000_00000;
		3090: oled_colour = 16'b00000_000000_00000;
		3091: oled_colour = 16'b00000_000000_00000;
		3092: oled_colour = 16'b00000_000000_00000;
		3093: oled_colour = 16'b00000_000000_00000;
		3094: oled_colour = 16'b00000_000000_00000;
		3095: oled_colour = 16'b00000_000000_00000;
		3096: oled_colour = 16'b00000_000000_00000;
		3097: oled_colour = 16'b00000_000000_00000;
		3098: oled_colour = 16'b00000_000000_00000;
		3099: oled_colour = 16'b00000_000000_00000;
		3100: oled_colour = 16'b00000_000000_00000;
		3101: oled_colour = 16'b00000_000000_00000;
		3102: oled_colour = 16'b00000_000000_00000;
		3103: oled_colour = 16'b00000_000000_00000;
		3104: oled_colour = 16'b00000_000000_00000;
		3105: oled_colour = 16'b00000_000000_00000;
		3106: oled_colour = 16'b00000_000000_00000;
		3107: oled_colour = 16'b00000_000000_00000;
		3108: oled_colour = 16'b00000_000000_00000;
		3109: oled_colour = 16'b00000_000000_00000;
		3110: oled_colour = 16'b00000_000000_00000;
		3111: oled_colour = 16'b00000_000000_00000;
		3112: oled_colour = 16'b00000_000000_00000;
		3113: oled_colour = 16'b11111_111111_11111; 
		3114: oled_colour = 16'b00000_000000_00000;
		3115: oled_colour = 16'b11101_111101_11101; 
		3116: oled_colour = 16'b10111_110001_10100; 
		3117: oled_colour = 16'b11001_101111_10011; 
		3118: oled_colour = 16'b11110_110111_10111; 
		3119: oled_colour = 16'b11001_110010_10110; 
		3120: oled_colour = 16'b10000_100111_01111; 
		3121: oled_colour = 16'b00101_010100_00010; 
		3122: oled_colour = 16'b10000_100001_01010; 
		3123: oled_colour = 16'b11010_110001_10101; 
		3124: oled_colour = 16'b11111_111111_11111; 
		3125: oled_colour = 16'b00000_000000_00000;
		3126: oled_colour = 16'b00000_000000_00000;
		3127: oled_colour = 16'b00000_000000_00000;
		3128: oled_colour = 16'b00000_000000_00000;
		3129: oled_colour = 16'b00000_000000_00000;
		3130: oled_colour = 16'b00000_000000_00000;
		3131: oled_colour = 16'b00000_000000_00000;
		3132: oled_colour = 16'b00000_000000_00000;
		3133: oled_colour = 16'b00000_000000_00000;
		3134: oled_colour = 16'b00000_000000_00000;
		3135: oled_colour = 16'b00000_000000_00000;
		3136: oled_colour = 16'b00000_000000_00000;
		3137: oled_colour = 16'b00000_000000_00000;
		3138: oled_colour = 16'b00000_000000_00000;
		3139: oled_colour = 16'b00000_000000_00000;
		3140: oled_colour = 16'b00000_000000_00000;
		3141: oled_colour = 16'b00000_000000_00000;
		3142: oled_colour = 16'b00000_000000_00000;
		3143: oled_colour = 16'b00000_000000_00000;
		3144: oled_colour = 16'b00000_000000_00000;
		3145: oled_colour = 16'b00000_000000_00000;
		3146: oled_colour = 16'b00000_000000_00000;
		3147: oled_colour = 16'b00000_000000_00000;
		3148: oled_colour = 16'b00000_000000_00000;
		3149: oled_colour = 16'b00000_000000_00000;
		3150: oled_colour = 16'b00000_000000_00000;
		3151: oled_colour = 16'b00000_000000_00000;
		3152: oled_colour = 16'b00000_000000_00000;
		3153: oled_colour = 16'b00000_000000_00000;
		3154: oled_colour = 16'b00000_000000_00000;
		3155: oled_colour = 16'b00000_000000_00000;
		3156: oled_colour = 16'b00000_000000_00000;
		3157: oled_colour = 16'b00000_000000_00000;
		3158: oled_colour = 16'b00000_000000_00000;
		3159: oled_colour = 16'b00000_000000_00000;
		3160: oled_colour = 16'b00000_000000_00000;
		3161: oled_colour = 16'b00000_000000_00000;
		3162: oled_colour = 16'b00000_000000_00000;
		3163: oled_colour = 16'b00000_000000_00000;
		3164: oled_colour = 16'b00000_000000_00000;
		3165: oled_colour = 16'b00000_000000_00000;
		3166: oled_colour = 16'b00000_000000_00000;
		3167: oled_colour = 16'b00000_000000_00000;
		3168: oled_colour = 16'b00000_000000_00000;
		3169: oled_colour = 16'b00000_000000_00000;
		3170: oled_colour = 16'b00000_000000_00000;
		3171: oled_colour = 16'b00000_000000_00000;
		3172: oled_colour = 16'b00000_000000_00000;
		3173: oled_colour = 16'b00000_000000_00000;
		3174: oled_colour = 16'b00000_000000_00000;
		3175: oled_colour = 16'b00000_000000_00000;
		3176: oled_colour = 16'b00000_000000_00000;
		3177: oled_colour = 16'b00000_000000_00000;
		3178: oled_colour = 16'b00000_000000_00000;
		3179: oled_colour = 16'b00000_000000_00000;
		3180: oled_colour = 16'b00000_000000_00000;
		3181: oled_colour = 16'b00000_000000_00000;
		3182: oled_colour = 16'b00000_000000_00000;
		3183: oled_colour = 16'b00000_000000_00000;
		3184: oled_colour = 16'b00000_000000_00000;
		3185: oled_colour = 16'b00000_000000_00000;
		3186: oled_colour = 16'b00000_000000_00000;
		3187: oled_colour = 16'b00000_000000_00000;
		3188: oled_colour = 16'b00000_000000_00000;
		3189: oled_colour = 16'b00000_000000_00000;
		3190: oled_colour = 16'b00000_000000_00000;
		3191: oled_colour = 16'b00000_000000_00000;
		3192: oled_colour = 16'b00000_000000_00000;
		3193: oled_colour = 16'b00000_000000_00000;
		3194: oled_colour = 16'b00000_000000_00000;
		3195: oled_colour = 16'b00000_000000_00000;
		3196: oled_colour = 16'b00000_000000_00000;
		3197: oled_colour = 16'b00000_000000_00000;
		3198: oled_colour = 16'b00000_000000_00000;
		3199: oled_colour = 16'b00000_000000_00000;
		3200: oled_colour = 16'b00000_000000_00000;
		3201: oled_colour = 16'b00000_000000_00000;
		3202: oled_colour = 16'b00000_000000_00000;
		3203: oled_colour = 16'b00000_000000_00000;
		3204: oled_colour = 16'b00000_000000_00000;
		3205: oled_colour = 16'b00000_000000_00000;
		3206: oled_colour = 16'b00000_000000_00000;
		3207: oled_colour = 16'b00000_000000_00000;
		3208: oled_colour = 16'b00000_000000_00000;
		3209: oled_colour = 16'b11111_111111_11111; 
		3210: oled_colour = 16'b00000_000000_00000;
		3211: oled_colour = 16'b11101_110111_11011; 
		3212: oled_colour = 16'b11100_101111_10100; 
		3213: oled_colour = 16'b11100_110000_10101; 
		3214: oled_colour = 16'b11101_101011_10010; 
		3215: oled_colour = 16'b11111_110100_10011; 
		3216: oled_colour = 16'b11001_101110_10010; 
		3217: oled_colour = 16'b00101_010110_00100; 
		3218: oled_colour = 16'b10111_101001_10001; 
		3219: oled_colour = 16'b11110_110101_11000; 
		3220: oled_colour = 16'b11110_111010_11101; 
		3221: oled_colour = 16'b11111_111111_11111; 
		3222: oled_colour = 16'b11111_111111_11111; 
		3223: oled_colour = 16'b00000_000000_00000;
		3224: oled_colour = 16'b00000_000000_00000;
		3225: oled_colour = 16'b00000_000000_00000;
		3226: oled_colour = 16'b00000_000000_00000;
		3227: oled_colour = 16'b00000_000000_00000;
		3228: oled_colour = 16'b00000_000000_00000;
		3229: oled_colour = 16'b00000_000000_00000;
		3230: oled_colour = 16'b00000_000000_00000;
		3231: oled_colour = 16'b00000_000000_00000;
		3232: oled_colour = 16'b00000_000000_00000;
		3233: oled_colour = 16'b00000_000000_00000;
		3234: oled_colour = 16'b00000_000000_00000;
		3235: oled_colour = 16'b00000_000000_00000;
		3236: oled_colour = 16'b00000_000000_00000;
		3237: oled_colour = 16'b00000_000000_00000;
		3238: oled_colour = 16'b00000_000000_00000;
		3239: oled_colour = 16'b00000_000000_00000;
		3240: oled_colour = 16'b00000_000000_00000;
		3241: oled_colour = 16'b00000_000000_00000;
		3242: oled_colour = 16'b00000_000000_00000;
		3243: oled_colour = 16'b00000_000000_00000;
		3244: oled_colour = 16'b00000_000000_00000;
		3245: oled_colour = 16'b00000_000000_00000;
		3246: oled_colour = 16'b00000_000000_00000;
		3247: oled_colour = 16'b00000_000000_00000;
		3248: oled_colour = 16'b00000_000000_00000;
		3249: oled_colour = 16'b00000_000000_00000;
		3250: oled_colour = 16'b00000_000000_00000;
		3251: oled_colour = 16'b00000_000000_00000;
		3252: oled_colour = 16'b00000_000000_00000;
		3253: oled_colour = 16'b00000_000000_00000;
		3254: oled_colour = 16'b00000_000000_00000;
		3255: oled_colour = 16'b00000_000000_00000;
		3256: oled_colour = 16'b00000_000000_00000;
		3257: oled_colour = 16'b00000_000000_00000;
		3258: oled_colour = 16'b00000_000000_00000;
		3259: oled_colour = 16'b00000_000000_00000;
		3260: oled_colour = 16'b00000_000000_00000;
		3261: oled_colour = 16'b00000_000000_00000;
		3262: oled_colour = 16'b00000_000000_00000;
		3263: oled_colour = 16'b00000_000000_00000;
		3264: oled_colour = 16'b00000_000000_00000;
		3265: oled_colour = 16'b00000_000000_00000;
		3266: oled_colour = 16'b00000_000000_00000;
		3267: oled_colour = 16'b00000_000000_00000;
		3268: oled_colour = 16'b00000_000000_00000;
		3269: oled_colour = 16'b00000_000000_00000;
		3270: oled_colour = 16'b00000_000000_00000;
		3271: oled_colour = 16'b00000_000000_00000;
		3272: oled_colour = 16'b00000_000000_00000;
		3273: oled_colour = 16'b00000_000000_00000;
		3274: oled_colour = 16'b00000_000000_00000;
		3275: oled_colour = 16'b00000_000000_00000;
		3276: oled_colour = 16'b00000_000000_00000;
		3277: oled_colour = 16'b00000_000000_00000;
		3278: oled_colour = 16'b00000_000000_00000;
		3279: oled_colour = 16'b00000_000000_00000;
		3280: oled_colour = 16'b00000_000000_00000;
		3281: oled_colour = 16'b00000_000000_00000;
		3282: oled_colour = 16'b00000_000000_00000;
		3283: oled_colour = 16'b00000_000000_00000;
		3284: oled_colour = 16'b00000_000000_00000;
		3285: oled_colour = 16'b00000_000000_00000;
		3286: oled_colour = 16'b00000_000000_00000;
		3287: oled_colour = 16'b00000_000000_00000;
		3288: oled_colour = 16'b00000_000000_00000;
		3289: oled_colour = 16'b00000_000000_00000;
		3290: oled_colour = 16'b00000_000000_00000;
		3291: oled_colour = 16'b00000_000000_00000;
		3292: oled_colour = 16'b00000_000000_00000;
		3293: oled_colour = 16'b00000_000000_00000;
		3294: oled_colour = 16'b00000_000000_00000;
		3295: oled_colour = 16'b00000_000000_00000;
		3296: oled_colour = 16'b00000_000000_00000;
		3297: oled_colour = 16'b00000_000000_00000;
		3298: oled_colour = 16'b00000_000000_00000;
		3299: oled_colour = 16'b00000_000000_00000;
		3300: oled_colour = 16'b00000_000000_00000;
		3301: oled_colour = 16'b00000_000000_00000;
		3302: oled_colour = 16'b00000_000000_00000;
		3303: oled_colour = 16'b00000_000000_00000;
		3304: oled_colour = 16'b00000_000000_00000;
		3305: oled_colour = 16'b11111_111111_11111; 
		3306: oled_colour = 16'b11111_111111_11111; 
		3307: oled_colour = 16'b11110_111001_11100; 
		3308: oled_colour = 16'b10010_101010_10001; 
		3309: oled_colour = 16'b10010_101111_10010; 
		3310: oled_colour = 16'b11011_110011_10010; 
		3311: oled_colour = 16'b11110_110100_10010; 
		3312: oled_colour = 16'b10110_110110_10010; 
		3313: oled_colour = 16'b01001_011100_01000; 
		3314: oled_colour = 16'b10110_110001_10010; 
		3315: oled_colour = 16'b11011_110101_10010; 
		3316: oled_colour = 16'b11100_101111_10101; 
		3317: oled_colour = 16'b00000_000000_00000;
		3318: oled_colour = 16'b11111_111111_11111; 
		3319: oled_colour = 16'b00000_000000_00000;
		3320: oled_colour = 16'b00000_000000_00000;
		3321: oled_colour = 16'b00000_000000_00000;
		3322: oled_colour = 16'b00000_000000_00000;
		3323: oled_colour = 16'b00000_000000_00000;
		3324: oled_colour = 16'b00000_000000_00000;
		3325: oled_colour = 16'b00000_000000_00000;
		3326: oled_colour = 16'b00000_000000_00000;
		3327: oled_colour = 16'b00000_000000_00000;
		3328: oled_colour = 16'b00000_000000_00000;
		3329: oled_colour = 16'b00000_000000_00000;
		3330: oled_colour = 16'b00000_000000_00000;
		3331: oled_colour = 16'b00000_000000_00000;
		3332: oled_colour = 16'b00000_000000_00000;
		3333: oled_colour = 16'b00000_000000_00000;
		3334: oled_colour = 16'b00000_000000_00000;
		3335: oled_colour = 16'b00000_000000_00000;
		3336: oled_colour = 16'b00000_000000_00000;
		3337: oled_colour = 16'b00000_000000_00000;
		3338: oled_colour = 16'b00000_000000_00000;
		3339: oled_colour = 16'b00000_000000_00000;
		3340: oled_colour = 16'b00000_000000_00000;
		3341: oled_colour = 16'b00000_000000_00000;
		3342: oled_colour = 16'b00000_000000_00000;
		3343: oled_colour = 16'b00000_000000_00000;
		3344: oled_colour = 16'b00000_000000_00000;
		3345: oled_colour = 16'b00000_000000_00000;
		3346: oled_colour = 16'b00000_000000_00000;
		3347: oled_colour = 16'b00000_000000_00000;
		3348: oled_colour = 16'b00000_000000_00000;
		3349: oled_colour = 16'b00000_000000_00000;
		3350: oled_colour = 16'b00000_000000_00000;
		3351: oled_colour = 16'b00000_000000_00000;
		3352: oled_colour = 16'b00000_000000_00000;
		3353: oled_colour = 16'b00000_000000_00000;
		3354: oled_colour = 16'b00000_000000_00000;
		3355: oled_colour = 16'b00000_000000_00000;
		3356: oled_colour = 16'b00000_000000_00000;
		3357: oled_colour = 16'b00000_000000_00000;
		3358: oled_colour = 16'b00000_000000_00000;
		3359: oled_colour = 16'b00000_000000_00000;
		3360: oled_colour = 16'b00000_000000_00000;
		3361: oled_colour = 16'b00000_000000_00000;
		3362: oled_colour = 16'b00000_000000_00000;
		3363: oled_colour = 16'b00000_000000_00000;
		3364: oled_colour = 16'b00000_000000_00000;
		3365: oled_colour = 16'b00000_000000_00000;
		3366: oled_colour = 16'b00000_000000_00000;
		3367: oled_colour = 16'b00000_000000_00000;
		3368: oled_colour = 16'b00000_000000_00000;
		3369: oled_colour = 16'b00000_000000_00000;
		3370: oled_colour = 16'b00000_000000_00000;
		3371: oled_colour = 16'b00000_000000_00000;
		3372: oled_colour = 16'b00000_000000_00000;
		3373: oled_colour = 16'b00000_000000_00000;
		3374: oled_colour = 16'b00000_000000_00000;
		3375: oled_colour = 16'b00000_000000_00000;
		3376: oled_colour = 16'b00000_000000_00000;
		3377: oled_colour = 16'b00000_000000_00000;
		3378: oled_colour = 16'b00000_000000_00000;
		3379: oled_colour = 16'b00000_000000_00000;
		3380: oled_colour = 16'b00000_000000_00000;
		3381: oled_colour = 16'b00000_000000_00000;
		3382: oled_colour = 16'b00000_000000_00000;
		3383: oled_colour = 16'b00000_000000_00000;
		3384: oled_colour = 16'b00000_000000_00000;
		3385: oled_colour = 16'b00000_000000_00000;
		3386: oled_colour = 16'b00000_000000_00000;
		3387: oled_colour = 16'b00000_000000_00000;
		3388: oled_colour = 16'b00000_000000_00000;
		3389: oled_colour = 16'b00000_000000_00000;
		3390: oled_colour = 16'b00000_000000_00000;
		3391: oled_colour = 16'b00000_000000_00000;
		3392: oled_colour = 16'b00000_000000_00000;
		3393: oled_colour = 16'b00000_000000_00000;
		3394: oled_colour = 16'b00000_000000_00000;
		3395: oled_colour = 16'b00000_000000_00000;
		3396: oled_colour = 16'b00000_000000_00000;
		3397: oled_colour = 16'b00000_000000_00000;
		3398: oled_colour = 16'b00000_000000_00000;
		3399: oled_colour = 16'b00000_000000_00000;
		3400: oled_colour = 16'b00000_000000_00000;
		3401: oled_colour = 16'b00000_000000_00000;
		3402: oled_colour = 16'b11111_111111_11111; 
		3403: oled_colour = 16'b00000_000000_00000;
		3404: oled_colour = 16'b11001_110110_11010; 
		3405: oled_colour = 16'b01100_100011_01011; 
		3406: oled_colour = 16'b10011_101011_01101; 
		3407: oled_colour = 16'b11100_110001_10011; 
		3408: oled_colour = 16'b11100_110100_10101; 
		3409: oled_colour = 16'b01100_100000_01011; 
		3410: oled_colour = 16'b10100_101101_10000; 
		3411: oled_colour = 16'b11111_111001_10111; 
		3412: oled_colour = 16'b11011_101111_10011; 
		3413: oled_colour = 16'b11111_111100_11110; 
		3414: oled_colour = 16'b00000_000000_00000;
		3415: oled_colour = 16'b11111_111111_11111; 
		3416: oled_colour = 16'b00000_000000_00000;
		3417: oled_colour = 16'b00000_000000_00000;
		3418: oled_colour = 16'b00000_000000_00000;
		3419: oled_colour = 16'b00000_000000_00000;
		3420: oled_colour = 16'b00000_000000_00000;
		3421: oled_colour = 16'b00000_000000_00000;
		3422: oled_colour = 16'b00000_000000_00000;
		3423: oled_colour = 16'b00000_000000_00000;
		3424: oled_colour = 16'b00000_000000_00000;
		3425: oled_colour = 16'b00000_000000_00000;
		3426: oled_colour = 16'b00000_000000_00000;
		3427: oled_colour = 16'b00000_000000_00000;
		3428: oled_colour = 16'b00000_000000_00000;
		3429: oled_colour = 16'b00000_000000_00000;
		3430: oled_colour = 16'b00000_000000_00000;
		3431: oled_colour = 16'b00000_000000_00000;
		3432: oled_colour = 16'b00000_000000_00000;
		3433: oled_colour = 16'b00000_000000_00000;
		3434: oled_colour = 16'b00000_000000_00000;
		3435: oled_colour = 16'b00000_000000_00000;
		3436: oled_colour = 16'b00000_000000_00000;
		3437: oled_colour = 16'b00000_000000_00000;
		3438: oled_colour = 16'b00000_000000_00000;
		3439: oled_colour = 16'b00000_000000_00000;
		3440: oled_colour = 16'b00000_000000_00000;
		3441: oled_colour = 16'b00000_000000_00000;
		3442: oled_colour = 16'b00000_000000_00000;
		3443: oled_colour = 16'b00000_000000_00000;
		3444: oled_colour = 16'b00000_000000_00000;
		3445: oled_colour = 16'b00000_000000_00000;
		3446: oled_colour = 16'b00000_000000_00000;
		3447: oled_colour = 16'b00000_000000_00000;
		3448: oled_colour = 16'b00000_000000_00000;
		3449: oled_colour = 16'b00000_000000_00000;
		3450: oled_colour = 16'b00000_000000_00000;
		3451: oled_colour = 16'b00000_000000_00000;
		3452: oled_colour = 16'b00000_000000_00000;
		3453: oled_colour = 16'b00000_000000_00000;
		3454: oled_colour = 16'b00000_000000_00000;
		3455: oled_colour = 16'b00000_000000_00000;
		3456: oled_colour = 16'b00000_000000_00000;
		3457: oled_colour = 16'b00000_000000_00000;
		3458: oled_colour = 16'b00000_000000_00000;
		3459: oled_colour = 16'b00000_000000_00000;
		3460: oled_colour = 16'b00000_000000_00000;
		3461: oled_colour = 16'b00000_000000_00000;
		3462: oled_colour = 16'b00000_000000_00000;
		3463: oled_colour = 16'b00000_000000_00000;
		3464: oled_colour = 16'b00000_000000_00000;
		3465: oled_colour = 16'b00000_000000_00000;
		3466: oled_colour = 16'b00000_000000_00000;
		3467: oled_colour = 16'b00000_000000_00000;
		3468: oled_colour = 16'b00000_000000_00000;
		3469: oled_colour = 16'b00000_000000_00000;
		3470: oled_colour = 16'b00000_000000_00000;
		3471: oled_colour = 16'b00000_000000_00000;
		3472: oled_colour = 16'b00000_000000_00000;
		3473: oled_colour = 16'b00000_000000_00000;
		3474: oled_colour = 16'b00000_000000_00000;
		3475: oled_colour = 16'b00000_000000_00000;
		3476: oled_colour = 16'b00000_000000_00000;
		3477: oled_colour = 16'b00000_000000_00000;
		3478: oled_colour = 16'b00000_000000_00000;
		3479: oled_colour = 16'b00000_000000_00000;
		3480: oled_colour = 16'b00000_000000_00000;
		3481: oled_colour = 16'b00000_000000_00000;
		3482: oled_colour = 16'b00000_000000_00000;
		3483: oled_colour = 16'b00000_000000_00000;
		3484: oled_colour = 16'b00000_000000_00000;
		3485: oled_colour = 16'b00000_000000_00000;
		3486: oled_colour = 16'b00000_000000_00000;
		3487: oled_colour = 16'b00000_000000_00000;
		3488: oled_colour = 16'b00000_000000_00000;
		3489: oled_colour = 16'b00000_000000_00000;
		3490: oled_colour = 16'b00000_000000_00000;
		3491: oled_colour = 16'b00000_000000_00000;
		3492: oled_colour = 16'b00000_000000_00000;
		3493: oled_colour = 16'b00000_000000_00000;
		3494: oled_colour = 16'b00000_000000_00000;
		3495: oled_colour = 16'b00000_000000_00000;
		3496: oled_colour = 16'b00000_000000_00000;
		3497: oled_colour = 16'b00000_000000_00000;
		3498: oled_colour = 16'b00000_000000_00000;
		3499: oled_colour = 16'b11111_111111_11111; 
		3500: oled_colour = 16'b00000_000000_00000;
		3501: oled_colour = 16'b10101_100100_01110; 
		3502: oled_colour = 16'b01100_011010_00111; 
		3503: oled_colour = 16'b10111_110011_10011; 
		3504: oled_colour = 16'b11000_111010_10110; 
		3505: oled_colour = 16'b01000_011101_01000; 
		3506: oled_colour = 16'b10000_101100_01110; 
		3507: oled_colour = 16'b11110_111100_11010; 
		3508: oled_colour = 16'b10100_100100_01101; 
		3509: oled_colour = 16'b11101_111000_11011; 
		3510: oled_colour = 16'b00000_000000_00000;
		3511: oled_colour = 16'b11111_111111_11111; 
		3512: oled_colour = 16'b00000_000000_00000;
		3513: oled_colour = 16'b00000_000000_00000;
		3514: oled_colour = 16'b00000_000000_00000;
		3515: oled_colour = 16'b00000_000000_00000;
		3516: oled_colour = 16'b00000_000000_00000;
		3517: oled_colour = 16'b00000_000000_00000;
		3518: oled_colour = 16'b00000_000000_00000;
		3519: oled_colour = 16'b00000_000000_00000;
		3520: oled_colour = 16'b00000_000000_00000;
		3521: oled_colour = 16'b00000_000000_00000;
		3522: oled_colour = 16'b00000_000000_00000;
		3523: oled_colour = 16'b00000_000000_00000;
		3524: oled_colour = 16'b00000_000000_00000;
		3525: oled_colour = 16'b00000_000000_00000;
		3526: oled_colour = 16'b00000_000000_00000;
		3527: oled_colour = 16'b00000_000000_00000;
		3528: oled_colour = 16'b00000_000000_00000;
		3529: oled_colour = 16'b00000_000000_00000;
		3530: oled_colour = 16'b00000_000000_00000;
		3531: oled_colour = 16'b00000_000000_00000;
		3532: oled_colour = 16'b00000_000000_00000;
		3533: oled_colour = 16'b00000_000000_00000;
		3534: oled_colour = 16'b00000_000000_00000;
		3535: oled_colour = 16'b00000_000000_00000;
		3536: oled_colour = 16'b00000_000000_00000;
		3537: oled_colour = 16'b00000_000000_00000;
		3538: oled_colour = 16'b00000_000000_00000;
		3539: oled_colour = 16'b00000_000000_00000;
		3540: oled_colour = 16'b00000_000000_00000;
		3541: oled_colour = 16'b00000_000000_00000;
		3542: oled_colour = 16'b00000_000000_00000;
		3543: oled_colour = 16'b00000_000000_00000;
		3544: oled_colour = 16'b00000_000000_00000;
		3545: oled_colour = 16'b00000_000000_00000;
		3546: oled_colour = 16'b00000_000000_00000;
		3547: oled_colour = 16'b00000_000000_00000;
		3548: oled_colour = 16'b00000_000000_00000;
		3549: oled_colour = 16'b00000_000000_00000;
		3550: oled_colour = 16'b00000_000000_00000;
		3551: oled_colour = 16'b00000_000000_00000;
		3552: oled_colour = 16'b00000_000000_00000;
		3553: oled_colour = 16'b00000_000000_00000;
		3554: oled_colour = 16'b00000_000000_00000;
		3555: oled_colour = 16'b00000_000000_00000;
		3556: oled_colour = 16'b00000_000000_00000;
		3557: oled_colour = 16'b00000_000000_00000;
		3558: oled_colour = 16'b00000_000000_00000;
		3559: oled_colour = 16'b00000_000000_00000;
		3560: oled_colour = 16'b00000_000000_00000;
		3561: oled_colour = 16'b00000_000000_00000;
		3562: oled_colour = 16'b00000_000000_00000;
		3563: oled_colour = 16'b00000_000000_00000;
		3564: oled_colour = 16'b00000_000000_00000;
		3565: oled_colour = 16'b00000_000000_00000;
		3566: oled_colour = 16'b00000_000000_00000;
		3567: oled_colour = 16'b00000_000000_00000;
		3568: oled_colour = 16'b00000_000000_00000;
		3569: oled_colour = 16'b00000_000000_00000;
		3570: oled_colour = 16'b00000_000000_00000;
		3571: oled_colour = 16'b00000_000000_00000;
		3572: oled_colour = 16'b00000_000000_00000;
		3573: oled_colour = 16'b00000_000000_00000;
		3574: oled_colour = 16'b00000_000000_00000;
		3575: oled_colour = 16'b00000_000000_00000;
		3576: oled_colour = 16'b00000_000000_00000;
		3577: oled_colour = 16'b00000_000000_00000;
		3578: oled_colour = 16'b00000_000000_00000;
		3579: oled_colour = 16'b00000_000000_00000;
		3580: oled_colour = 16'b00000_000000_00000;
		3581: oled_colour = 16'b00000_000000_00000;
		3582: oled_colour = 16'b00000_000000_00000;
		3583: oled_colour = 16'b00000_000000_00000;
		3584: oled_colour = 16'b00000_000000_00000;
		3585: oled_colour = 16'b00000_000000_00000;
		3586: oled_colour = 16'b00000_000000_00000;
		3587: oled_colour = 16'b00000_000000_00000;
		3588: oled_colour = 16'b00000_000000_00000;
		3589: oled_colour = 16'b00000_000000_00000;
		3590: oled_colour = 16'b00000_000000_00000;
		3591: oled_colour = 16'b00000_000000_00000;
		3592: oled_colour = 16'b00000_000000_00000;
		3593: oled_colour = 16'b00000_000000_00000;
		3594: oled_colour = 16'b11111_111111_11111; 
		3595: oled_colour = 16'b00000_000000_00000;
		3596: oled_colour = 16'b11110_111100_11110; 
		3597: oled_colour = 16'b10110_100111_01110; 
		3598: oled_colour = 16'b11000_101101_10010; 
		3599: oled_colour = 16'b10101_110011_10101; 
		3600: oled_colour = 16'b10111_110010_10011; 
		3601: oled_colour = 16'b10000_011010_01000; 
		3602: oled_colour = 16'b01111_100111_10000; 
		3603: oled_colour = 16'b10011_101110_10000; 
		3604: oled_colour = 16'b10110_101011_10010; 
		3605: oled_colour = 16'b11111_111110_11111; 
		3606: oled_colour = 16'b11111_111111_11111; 
		3607: oled_colour = 16'b00000_000000_00000;
		3608: oled_colour = 16'b00000_000000_00000;
		3609: oled_colour = 16'b00000_000000_00000;
		3610: oled_colour = 16'b00000_000000_00000;
		3611: oled_colour = 16'b00000_000000_00000;
		3612: oled_colour = 16'b00000_000000_00000;
		3613: oled_colour = 16'b00000_000000_00000;
		3614: oled_colour = 16'b00000_000000_00000;
		3615: oled_colour = 16'b00000_000000_00000;
		3616: oled_colour = 16'b00000_000000_00000;
		3617: oled_colour = 16'b00000_000000_00000;
		3618: oled_colour = 16'b00000_000000_00000;
		3619: oled_colour = 16'b00000_000000_00000;
		3620: oled_colour = 16'b00000_000000_00000;
		3621: oled_colour = 16'b00000_000000_00000;
		3622: oled_colour = 16'b00000_000000_00000;
		3623: oled_colour = 16'b00000_000000_00000;
		3624: oled_colour = 16'b00000_000000_00000;
		3625: oled_colour = 16'b00000_000000_00000;
		3626: oled_colour = 16'b00000_000000_00000;
		3627: oled_colour = 16'b00000_000000_00000;
		3628: oled_colour = 16'b00000_000000_00000;
		3629: oled_colour = 16'b00000_000000_00000;
		3630: oled_colour = 16'b00000_000000_00000;
		3631: oled_colour = 16'b00000_000000_00000;
		3632: oled_colour = 16'b00000_000000_00000;
		3633: oled_colour = 16'b00000_000000_00000;
		3634: oled_colour = 16'b00000_000000_00000;
		3635: oled_colour = 16'b00000_000000_00000;
		3636: oled_colour = 16'b00000_000000_00000;
		3637: oled_colour = 16'b00000_000000_00000;
		3638: oled_colour = 16'b00000_000000_00000;
		3639: oled_colour = 16'b00000_000000_00000;
		3640: oled_colour = 16'b00000_000000_00000;
		3641: oled_colour = 16'b00000_000000_00000;
		3642: oled_colour = 16'b00000_000000_00000;
		3643: oled_colour = 16'b00000_000000_00000;
		3644: oled_colour = 16'b00000_000000_00000;
		3645: oled_colour = 16'b00000_000000_00000;
		3646: oled_colour = 16'b00000_000000_00000;
		3647: oled_colour = 16'b00000_000000_00000;
		3648: oled_colour = 16'b00000_000000_00000;
		3649: oled_colour = 16'b00000_000000_00000;
		3650: oled_colour = 16'b00000_000000_00000;
		3651: oled_colour = 16'b00000_000000_00000;
		3652: oled_colour = 16'b00000_000000_00000;
		3653: oled_colour = 16'b00000_000000_00000;
		3654: oled_colour = 16'b00000_000000_00000;
		3655: oled_colour = 16'b00000_000000_00000;
		3656: oled_colour = 16'b00000_000000_00000;
		3657: oled_colour = 16'b00000_000000_00000;
		3658: oled_colour = 16'b00000_000000_00000;
		3659: oled_colour = 16'b00000_000000_00000;
		3660: oled_colour = 16'b00000_000000_00000;
		3661: oled_colour = 16'b00000_000000_00000;
		3662: oled_colour = 16'b00000_000000_00000;
		3663: oled_colour = 16'b00000_000000_00000;
		3664: oled_colour = 16'b00000_000000_00000;
		3665: oled_colour = 16'b00000_000000_00000;
		3666: oled_colour = 16'b00000_000000_00000;
		3667: oled_colour = 16'b00000_000000_00000;
		3668: oled_colour = 16'b00000_000000_00000;
		3669: oled_colour = 16'b00000_000000_00000;
		3670: oled_colour = 16'b00000_000000_00000;
		3671: oled_colour = 16'b00000_000000_00000;
		3672: oled_colour = 16'b00000_000000_00000;
		3673: oled_colour = 16'b00000_000000_00000;
		3674: oled_colour = 16'b00000_000000_00000;
		3675: oled_colour = 16'b00000_000000_00000;
		3676: oled_colour = 16'b00000_000000_00000;
		3677: oled_colour = 16'b00000_000000_00000;
		3678: oled_colour = 16'b00000_000000_00000;
		3679: oled_colour = 16'b00000_000000_00000;
		3680: oled_colour = 16'b00000_000000_00000;
		3681: oled_colour = 16'b00000_000000_00000;
		3682: oled_colour = 16'b00000_000000_00000;
		3683: oled_colour = 16'b00000_000000_00000;
		3684: oled_colour = 16'b00000_000000_00000;
		3685: oled_colour = 16'b00000_000000_00000;
		3686: oled_colour = 16'b00000_000000_00000;
		3687: oled_colour = 16'b00000_000000_00000;
		3688: oled_colour = 16'b00000_000000_00000;
		3689: oled_colour = 16'b00000_000000_00000;
		3690: oled_colour = 16'b11111_111111_11111; 
		3691: oled_colour = 16'b00000_000000_00000;
		3692: oled_colour = 16'b11111_111100_11110; 
		3693: oled_colour = 16'b01110_011110_01001; 
		3694: oled_colour = 16'b10100_110001_10011; 
		3695: oled_colour = 16'b11001_110000_10100; 
		3696: oled_colour = 16'b10001_100000_01011; 
		3697: oled_colour = 16'b01011_010110_00101; 
		3698: oled_colour = 16'b10001_100000_01011; 
		3699: oled_colour = 16'b11010_110011_10111; 
		3700: oled_colour = 16'b00000_000000_00000;
		3701: oled_colour = 16'b00000_000000_00000;
		3702: oled_colour = 16'b00000_000000_00000;
		3703: oled_colour = 16'b00000_000000_00000;
		3704: oled_colour = 16'b00000_000000_00000;
		3705: oled_colour = 16'b00000_000000_00000;
		3706: oled_colour = 16'b00000_000000_00000;
		3707: oled_colour = 16'b00000_000000_00000;
		3708: oled_colour = 16'b00000_000000_00000;
		3709: oled_colour = 16'b00000_000000_00000;
		3710: oled_colour = 16'b00000_000000_00000;
		3711: oled_colour = 16'b00000_000000_00000;
		3712: oled_colour = 16'b00000_000000_00000;
		3713: oled_colour = 16'b00000_000000_00000;
		3714: oled_colour = 16'b00000_000000_00000;
		3715: oled_colour = 16'b00000_000000_00000;
		3716: oled_colour = 16'b00000_000000_00000;
		3717: oled_colour = 16'b00000_000000_00000;
		3718: oled_colour = 16'b00000_000000_00000;
		3719: oled_colour = 16'b00000_000000_00000;
		3720: oled_colour = 16'b00000_000000_00000;
		3721: oled_colour = 16'b00000_000000_00000;
		3722: oled_colour = 16'b00000_000000_00000;
		3723: oled_colour = 16'b00000_000000_00000;
		3724: oled_colour = 16'b00000_000000_00000;
		3725: oled_colour = 16'b00000_000000_00000;
		3726: oled_colour = 16'b00000_000000_00000;
		3727: oled_colour = 16'b00000_000000_00000;
		3728: oled_colour = 16'b00000_000000_00000;
		3729: oled_colour = 16'b00000_000000_00000;
		3730: oled_colour = 16'b00000_000000_00000;
		3731: oled_colour = 16'b00000_000000_00000;
		3732: oled_colour = 16'b00000_000000_00000;
		3733: oled_colour = 16'b00000_000000_00000;
		3734: oled_colour = 16'b00000_000000_00000;
		3735: oled_colour = 16'b00000_000000_00000;
		3736: oled_colour = 16'b00000_000000_00000;
		3737: oled_colour = 16'b00000_000000_00000;
		3738: oled_colour = 16'b00000_000000_00000;
		3739: oled_colour = 16'b00000_000000_00000;
		3740: oled_colour = 16'b00000_000000_00000;
		3741: oled_colour = 16'b00000_000000_00000;
		3742: oled_colour = 16'b00000_000000_00000;
		3743: oled_colour = 16'b00000_000000_00000;
		3744: oled_colour = 16'b00000_000000_00000;
		3745: oled_colour = 16'b00000_000000_00000;
		3746: oled_colour = 16'b00000_000000_00000;
		3747: oled_colour = 16'b00000_000000_00000;
		3748: oled_colour = 16'b00000_000000_00000;
		3749: oled_colour = 16'b00000_000000_00000;
		3750: oled_colour = 16'b00000_000000_00000;
		3751: oled_colour = 16'b00000_000000_00000;
		3752: oled_colour = 16'b00000_000000_00000;
		3753: oled_colour = 16'b00000_000000_00000;
		3754: oled_colour = 16'b00000_000000_00000;
		3755: oled_colour = 16'b00000_000000_00000;
		3756: oled_colour = 16'b00000_000000_00000;
		3757: oled_colour = 16'b00000_000000_00000;
		3758: oled_colour = 16'b00000_000000_00000;
		3759: oled_colour = 16'b00000_000000_00000;
		3760: oled_colour = 16'b00000_000000_00000;
		3761: oled_colour = 16'b00000_000000_00000;
		3762: oled_colour = 16'b00000_000000_00000;
		3763: oled_colour = 16'b00000_000000_00000;
		3764: oled_colour = 16'b00000_000000_00000;
		3765: oled_colour = 16'b00000_000000_00000;
		3766: oled_colour = 16'b00000_000000_00000;
		3767: oled_colour = 16'b00000_000000_00000;
		3768: oled_colour = 16'b00000_000000_00000;
		3769: oled_colour = 16'b00000_000000_00000;
		3770: oled_colour = 16'b00000_000000_00000;
		3771: oled_colour = 16'b00000_000000_00000;
		3772: oled_colour = 16'b00000_000000_00000;
		3773: oled_colour = 16'b00000_000000_00000;
		3774: oled_colour = 16'b00000_000000_00000;
		3775: oled_colour = 16'b00000_000000_00000;
		3776: oled_colour = 16'b00000_000000_00000;
		3777: oled_colour = 16'b00000_000000_00000;
		3778: oled_colour = 16'b00000_000000_00000;
		3779: oled_colour = 16'b00000_000000_00000;
		3780: oled_colour = 16'b00000_000000_00000;
		3781: oled_colour = 16'b00000_000000_00000;
		3782: oled_colour = 16'b00000_000000_00000;
		3783: oled_colour = 16'b00000_000000_00000;
		3784: oled_colour = 16'b00000_000000_00000;
		3785: oled_colour = 16'b00000_000000_00000;
		3786: oled_colour = 16'b00000_000000_00000;
		3787: oled_colour = 16'b11111_111111_11111; 
		3788: oled_colour = 16'b00000_000000_00000;
		3789: oled_colour = 16'b10101_101001_10001; 
		3790: oled_colour = 16'b01010_010110_00100; 
		3791: oled_colour = 16'b01011_011101_00111; 
		3792: oled_colour = 16'b01010_010011_00010; 
		3793: oled_colour = 16'b01111_010110_00101; 
		3794: oled_colour = 16'b10110_101010_10010; 
		3795: oled_colour = 16'b00000_000000_00000;
		3796: oled_colour = 16'b11111_111111_11111; 
		3797: oled_colour = 16'b11111_111111_11111; 
		3798: oled_colour = 16'b00000_000000_00000;
		3799: oled_colour = 16'b00000_000000_00000;
		3800: oled_colour = 16'b00000_000000_00000;
		3801: oled_colour = 16'b00000_000000_00000;
		3802: oled_colour = 16'b00000_000000_00000;
		3803: oled_colour = 16'b00000_000000_00000;
		3804: oled_colour = 16'b00000_000000_00000;
		3805: oled_colour = 16'b00000_000000_00000;
		3806: oled_colour = 16'b00000_000000_00000;
		3807: oled_colour = 16'b00000_000000_00000;
		3808: oled_colour = 16'b00000_000000_00000;
		3809: oled_colour = 16'b00000_000000_00000;
		3810: oled_colour = 16'b00000_000000_00000;
		3811: oled_colour = 16'b00000_000000_00000;
		3812: oled_colour = 16'b00000_000000_00000;
		3813: oled_colour = 16'b00000_000000_00000;
		3814: oled_colour = 16'b00000_000000_00000;
		3815: oled_colour = 16'b00000_000000_00000;
		3816: oled_colour = 16'b00000_000000_00000;
		3817: oled_colour = 16'b00000_000000_00000;
		3818: oled_colour = 16'b00000_000000_00000;
		3819: oled_colour = 16'b00000_000000_00000;
		3820: oled_colour = 16'b00000_000000_00000;
		3821: oled_colour = 16'b00000_000000_00000;
		3822: oled_colour = 16'b00000_000000_00000;
		3823: oled_colour = 16'b00000_000000_00000;
		3824: oled_colour = 16'b00000_000000_00000;
		3825: oled_colour = 16'b00000_000000_00000;
		3826: oled_colour = 16'b00000_000000_00000;
		3827: oled_colour = 16'b00000_000000_00000;
		3828: oled_colour = 16'b00000_000000_00000;
		3829: oled_colour = 16'b00000_000000_00000;
		3830: oled_colour = 16'b00000_000000_00000;
		3831: oled_colour = 16'b00000_000000_00000;
		3832: oled_colour = 16'b00000_000000_00000;
		3833: oled_colour = 16'b00000_000000_00000;
		3834: oled_colour = 16'b00000_000000_00000;
		3835: oled_colour = 16'b00000_000000_00000;
		3836: oled_colour = 16'b00000_000000_00000;
		3837: oled_colour = 16'b00000_000000_00000;
		3838: oled_colour = 16'b00000_000000_00000;
		3839: oled_colour = 16'b00000_000000_00000;
		3840: oled_colour = 16'b00000_000000_00000;
		3841: oled_colour = 16'b00000_000000_00000;
		3842: oled_colour = 16'b00000_000000_00000;
		3843: oled_colour = 16'b00000_000000_00000;
		3844: oled_colour = 16'b00000_000000_00000;
		3845: oled_colour = 16'b00000_000000_00000;
		3846: oled_colour = 16'b00000_000000_00000;
		3847: oled_colour = 16'b00000_000000_00000;
		3848: oled_colour = 16'b00000_000000_00000;
		3849: oled_colour = 16'b00000_000000_00000;
		3850: oled_colour = 16'b00000_000000_00000;
		3851: oled_colour = 16'b00000_000000_00000;
		3852: oled_colour = 16'b00000_000000_00000;
		3853: oled_colour = 16'b00000_000000_00000;
		3854: oled_colour = 16'b00000_000000_00000;
		3855: oled_colour = 16'b00000_000000_00000;
		3856: oled_colour = 16'b00000_000000_00000;
		3857: oled_colour = 16'b00000_000000_00000;
		3858: oled_colour = 16'b00000_000000_00000;
		3859: oled_colour = 16'b00000_000000_00000;
		3860: oled_colour = 16'b00000_000000_00000;
		3861: oled_colour = 16'b00000_000000_00000;
		3862: oled_colour = 16'b00000_000000_00000;
		3863: oled_colour = 16'b00000_000000_00000;
		3864: oled_colour = 16'b00000_000000_00000;
		3865: oled_colour = 16'b00000_000000_00000;
		3866: oled_colour = 16'b00000_000000_00000;
		3867: oled_colour = 16'b00000_000000_00000;
		3868: oled_colour = 16'b00000_000000_00000;
		3869: oled_colour = 16'b00000_000000_00000;
		3870: oled_colour = 16'b00000_000000_00000;
		3871: oled_colour = 16'b00000_000000_00000;
		3872: oled_colour = 16'b00000_000000_00000;
		3873: oled_colour = 16'b00000_000000_00000;
		3874: oled_colour = 16'b00000_000000_00000;
		3875: oled_colour = 16'b00000_000000_00000;
		3876: oled_colour = 16'b00000_000000_00000;
		3877: oled_colour = 16'b00000_000000_00000;
		3878: oled_colour = 16'b00000_000000_00000;
		3879: oled_colour = 16'b00000_000000_00000;
		3880: oled_colour = 16'b00000_000000_00000;
		3881: oled_colour = 16'b00000_000000_00000;
		3882: oled_colour = 16'b00000_000000_00000;
		3883: oled_colour = 16'b11111_111111_11111; 
		3884: oled_colour = 16'b00000_000000_00000;
		3885: oled_colour = 16'b10111_101011_10011; 
		3886: oled_colour = 16'b10001_010110_00101; 
		3887: oled_colour = 16'b10001_010110_00101; 
		3888: oled_colour = 16'b01110_010001_00010; 
		3889: oled_colour = 16'b10110_100000_01100; 
		3890: oled_colour = 16'b11111_111111_11111; 
		3891: oled_colour = 16'b11111_111111_11111; 
		3892: oled_colour = 16'b11111_111111_11111; 
		3893: oled_colour = 16'b00000_000000_00000;
		3894: oled_colour = 16'b00000_000000_00000;
		3895: oled_colour = 16'b00000_000000_00000;
		3896: oled_colour = 16'b00000_000000_00000;
		3897: oled_colour = 16'b00000_000000_00000;
		3898: oled_colour = 16'b00000_000000_00000;
		3899: oled_colour = 16'b00000_000000_00000;
		3900: oled_colour = 16'b00000_000000_00000;
		3901: oled_colour = 16'b00000_000000_00000;
		3902: oled_colour = 16'b00000_000000_00000;
		3903: oled_colour = 16'b00000_000000_00000;
		3904: oled_colour = 16'b00000_000000_00000;
		3905: oled_colour = 16'b00000_000000_00000;
		3906: oled_colour = 16'b00000_000000_00000;
		3907: oled_colour = 16'b00000_000000_00000;
		3908: oled_colour = 16'b00000_000000_00000;
		3909: oled_colour = 16'b00000_000000_00000;
		3910: oled_colour = 16'b00000_000000_00000;
		3911: oled_colour = 16'b00000_000000_00000;
		3912: oled_colour = 16'b00000_000000_00000;
		3913: oled_colour = 16'b00000_000000_00000;
		3914: oled_colour = 16'b00000_000000_00000;
		3915: oled_colour = 16'b00000_000000_00000;
		3916: oled_colour = 16'b00000_000000_00000;
		3917: oled_colour = 16'b00000_000000_00000;
		3918: oled_colour = 16'b00000_000000_00000;
		3919: oled_colour = 16'b00000_000000_00000;
		3920: oled_colour = 16'b00000_000000_00000;
		3921: oled_colour = 16'b00000_000000_00000;
		3922: oled_colour = 16'b00000_000000_00000;
		3923: oled_colour = 16'b00000_000000_00000;
		3924: oled_colour = 16'b00000_000000_00000;
		3925: oled_colour = 16'b00000_000000_00000;
		3926: oled_colour = 16'b00000_000000_00000;
		3927: oled_colour = 16'b00000_000000_00000;
		3928: oled_colour = 16'b00000_000000_00000;
		3929: oled_colour = 16'b00000_000000_00000;
		3930: oled_colour = 16'b00000_000000_00000;
		3931: oled_colour = 16'b00000_000000_00000;
		3932: oled_colour = 16'b00000_000000_00000;
		3933: oled_colour = 16'b00000_000000_00000;
		3934: oled_colour = 16'b00000_000000_00000;
		3935: oled_colour = 16'b00000_000000_00000;
		3936: oled_colour = 16'b00000_000000_00000;
		3937: oled_colour = 16'b00000_000000_00000;
		3938: oled_colour = 16'b00000_000000_00000;
		3939: oled_colour = 16'b00000_000000_00000;
		3940: oled_colour = 16'b00000_000000_00000;
		3941: oled_colour = 16'b00000_000000_00000;
		3942: oled_colour = 16'b00000_000000_00000;
		3943: oled_colour = 16'b00000_000000_00000;
		3944: oled_colour = 16'b00000_000000_00000;
		3945: oled_colour = 16'b00000_000000_00000;
		3946: oled_colour = 16'b00000_000000_00000;
		3947: oled_colour = 16'b00000_000000_00000;
		3948: oled_colour = 16'b00000_000000_00000;
		3949: oled_colour = 16'b00000_000000_00000;
		3950: oled_colour = 16'b00000_000000_00000;
		3951: oled_colour = 16'b00000_000000_00000;
		3952: oled_colour = 16'b00000_000000_00000;
		3953: oled_colour = 16'b00000_000000_00000;
		3954: oled_colour = 16'b00000_000000_00000;
		3955: oled_colour = 16'b00000_000000_00000;
		3956: oled_colour = 16'b00000_000000_00000;
		3957: oled_colour = 16'b00000_000000_00000;
		3958: oled_colour = 16'b00000_000000_00000;
		3959: oled_colour = 16'b00000_000000_00000;
		3960: oled_colour = 16'b00000_000000_00000;
		3961: oled_colour = 16'b00000_000000_00000;
		3962: oled_colour = 16'b00000_000000_00000;
		3963: oled_colour = 16'b00000_000000_00000;
		3964: oled_colour = 16'b00000_000000_00000;
		3965: oled_colour = 16'b00000_000000_00000;
		3966: oled_colour = 16'b00000_000000_00000;
		3967: oled_colour = 16'b00000_000000_00000;
		3968: oled_colour = 16'b00000_000000_00000;
		3969: oled_colour = 16'b00000_000000_00000;
		3970: oled_colour = 16'b00000_000000_00000;
		3971: oled_colour = 16'b00000_000000_00000;
		3972: oled_colour = 16'b00000_000000_00000;
		3973: oled_colour = 16'b00000_000000_00000;
		3974: oled_colour = 16'b00000_000000_00000;
		3975: oled_colour = 16'b00000_000000_00000;
		3976: oled_colour = 16'b00000_000000_00000;
		3977: oled_colour = 16'b00000_000000_00000;
		3978: oled_colour = 16'b00000_000000_00000;
		3979: oled_colour = 16'b11111_111111_11111; 
		3980: oled_colour = 16'b00000_000000_00000;
		3981: oled_colour = 16'b10111_101010_10010; 
		3982: oled_colour = 16'b10001_010110_00101; 
		3983: oled_colour = 16'b01111_010101_00100; 
		3984: oled_colour = 16'b01101_010001_00010; 
		3985: oled_colour = 16'b10100_011101_01010; 
		3986: oled_colour = 16'b11111_111110_11111; 
		3987: oled_colour = 16'b00000_000000_00000;
		3988: oled_colour = 16'b11111_111111_11111; 
		3989: oled_colour = 16'b00000_000000_00000;
		3990: oled_colour = 16'b00000_000000_00000;
		3991: oled_colour = 16'b00000_000000_00000;
		3992: oled_colour = 16'b00000_000000_00000;
		3993: oled_colour = 16'b00000_000000_00000;
		3994: oled_colour = 16'b00000_000000_00000;
		3995: oled_colour = 16'b00000_000000_00000;
		3996: oled_colour = 16'b00000_000000_00000;
		3997: oled_colour = 16'b00000_000000_00000;
		3998: oled_colour = 16'b00000_000000_00000;
		3999: oled_colour = 16'b00000_000000_00000;
		4000: oled_colour = 16'b00000_000000_00000;
		4001: oled_colour = 16'b00000_000000_00000;
		4002: oled_colour = 16'b00000_000000_00000;
		4003: oled_colour = 16'b00000_000000_00000;
		4004: oled_colour = 16'b00000_000000_00000;
		4005: oled_colour = 16'b00000_000000_00000;
		4006: oled_colour = 16'b00000_000000_00000;
		4007: oled_colour = 16'b00000_000000_00000;
		4008: oled_colour = 16'b00000_000000_00000;
		4009: oled_colour = 16'b00000_000000_00000;
		4010: oled_colour = 16'b00000_000000_00000;
		4011: oled_colour = 16'b00000_000000_00000;
		4012: oled_colour = 16'b00000_000000_00000;
		4013: oled_colour = 16'b00000_000000_00000;
		4014: oled_colour = 16'b00000_000000_00000;
		4015: oled_colour = 16'b00000_000000_00000;
		4016: oled_colour = 16'b00000_000000_00000;
		4017: oled_colour = 16'b00000_000000_00000;
		4018: oled_colour = 16'b00000_000000_00000;
		4019: oled_colour = 16'b00000_000000_00000;
		4020: oled_colour = 16'b00000_000000_00000;
		4021: oled_colour = 16'b00000_000000_00000;
		4022: oled_colour = 16'b00000_000000_00000;
		4023: oled_colour = 16'b00000_000000_00000;
		4024: oled_colour = 16'b00000_000000_00000;
		4025: oled_colour = 16'b00000_000000_00000;
		4026: oled_colour = 16'b00000_000000_00000;
		4027: oled_colour = 16'b00000_000000_00000;
		4028: oled_colour = 16'b00000_000000_00000;
		4029: oled_colour = 16'b00000_000000_00000;
		4030: oled_colour = 16'b00000_000000_00000;
		4031: oled_colour = 16'b00000_000000_00000;
		4032: oled_colour = 16'b00000_000000_00000;
		4033: oled_colour = 16'b00000_000000_00000;
		4034: oled_colour = 16'b00000_000000_00000;
		4035: oled_colour = 16'b00000_000000_00000;
		4036: oled_colour = 16'b00000_000000_00000;
		4037: oled_colour = 16'b00000_000000_00000;
		4038: oled_colour = 16'b00000_000000_00000;
		4039: oled_colour = 16'b00000_000000_00000;
		4040: oled_colour = 16'b00000_000000_00000;
		4041: oled_colour = 16'b00000_000000_00000;
		4042: oled_colour = 16'b00000_000000_00000;
		4043: oled_colour = 16'b00000_000000_00000;
		4044: oled_colour = 16'b00000_000000_00000;
		4045: oled_colour = 16'b00000_000000_00000;
		4046: oled_colour = 16'b00000_000000_00000;
		4047: oled_colour = 16'b00000_000000_00000;
		4048: oled_colour = 16'b00000_000000_00000;
		4049: oled_colour = 16'b00000_000000_00000;
		4050: oled_colour = 16'b00000_000000_00000;
		4051: oled_colour = 16'b00000_000000_00000;
		4052: oled_colour = 16'b00000_000000_00000;
		4053: oled_colour = 16'b00000_000000_00000;
		4054: oled_colour = 16'b00000_000000_00000;
		4055: oled_colour = 16'b00000_000000_00000;
		4056: oled_colour = 16'b00000_000000_00000;
		4057: oled_colour = 16'b00000_000000_00000;
		4058: oled_colour = 16'b00000_000000_00000;
		4059: oled_colour = 16'b00000_000000_00000;
		4060: oled_colour = 16'b00000_000000_00000;
		4061: oled_colour = 16'b00000_000000_00000;
		4062: oled_colour = 16'b00000_000000_00000;
		4063: oled_colour = 16'b00000_000000_00000;
		4064: oled_colour = 16'b00000_000000_00000;
		4065: oled_colour = 16'b00000_000000_00000;
		4066: oled_colour = 16'b00000_000000_00000;
		4067: oled_colour = 16'b00000_000000_00000;
		4068: oled_colour = 16'b00000_000000_00000;
		4069: oled_colour = 16'b00000_000000_00000;
		4070: oled_colour = 16'b00000_000000_00000;
		4071: oled_colour = 16'b00000_000000_00000;
		4072: oled_colour = 16'b00000_000000_00000;
		4073: oled_colour = 16'b00000_000000_00000;
		4074: oled_colour = 16'b00000_000000_00000;
		4075: oled_colour = 16'b11111_111111_11111; 
		4076: oled_colour = 16'b00000_000000_00000;
		4077: oled_colour = 16'b10111_101011_10011; 
		4078: oled_colour = 16'b10010_011000_00110; 
		4079: oled_colour = 16'b01111_010100_00100; 
		4080: oled_colour = 16'b10100_011101_01001; 
		4081: oled_colour = 16'b11010_100111_01111; 
		4082: oled_colour = 16'b11100_110011_11000; 
		4083: oled_colour = 16'b00000_000000_00000;
		4084: oled_colour = 16'b11111_111111_11111; 
		4085: oled_colour = 16'b00000_000000_00000;
		4086: oled_colour = 16'b00000_000000_00000;
		4087: oled_colour = 16'b00000_000000_00000;
		4088: oled_colour = 16'b00000_000000_00000;
		4089: oled_colour = 16'b00000_000000_00000;
		4090: oled_colour = 16'b00000_000000_00000;
		4091: oled_colour = 16'b00000_000000_00000;
		4092: oled_colour = 16'b00000_000000_00000;
		4093: oled_colour = 16'b00000_000000_00000;
		4094: oled_colour = 16'b00000_000000_00000;
		4095: oled_colour = 16'b00000_000000_00000;
		4096: oled_colour = 16'b00000_000000_00000;
		4097: oled_colour = 16'b00000_000000_00000;
		4098: oled_colour = 16'b00000_000000_00000;
		4099: oled_colour = 16'b00000_000000_00000;
		4100: oled_colour = 16'b00000_000000_00000;
		4101: oled_colour = 16'b00000_000000_00000;
		4102: oled_colour = 16'b00000_000000_00000;
		4103: oled_colour = 16'b00000_000000_00000;
		4104: oled_colour = 16'b00000_000000_00000;
		4105: oled_colour = 16'b00000_000000_00000;
		4106: oled_colour = 16'b00000_000000_00000;
		4107: oled_colour = 16'b00000_000000_00000;
		4108: oled_colour = 16'b00000_000000_00000;
		4109: oled_colour = 16'b00000_000000_00000;
		4110: oled_colour = 16'b00000_000000_00000;
		4111: oled_colour = 16'b00000_000000_00000;
		4112: oled_colour = 16'b00000_000000_00000;
		4113: oled_colour = 16'b00000_000000_00000;
		4114: oled_colour = 16'b00000_000000_00000;
		4115: oled_colour = 16'b00000_000000_00000;
		4116: oled_colour = 16'b00000_000000_00000;
		4117: oled_colour = 16'b00000_000000_00000;
		4118: oled_colour = 16'b00000_000000_00000;
		4119: oled_colour = 16'b00000_000000_00000;
		4120: oled_colour = 16'b00000_000000_00000;
		4121: oled_colour = 16'b00000_000000_00000;
		4122: oled_colour = 16'b00000_000000_00000;
		4123: oled_colour = 16'b00000_000000_00000;
		4124: oled_colour = 16'b00000_000000_00000;
		4125: oled_colour = 16'b00000_000000_00000;
		4126: oled_colour = 16'b00000_000000_00000;
		4127: oled_colour = 16'b00000_000000_00000;
		4128: oled_colour = 16'b00000_000000_00000;
		4129: oled_colour = 16'b00000_000000_00000;
		4130: oled_colour = 16'b00000_000000_00000;
		4131: oled_colour = 16'b00000_000000_00000;
		4132: oled_colour = 16'b00000_000000_00000;
		4133: oled_colour = 16'b00000_000000_00000;
		4134: oled_colour = 16'b00000_000000_00000;
		4135: oled_colour = 16'b00000_000000_00000;
		4136: oled_colour = 16'b00000_000000_00000;
		4137: oled_colour = 16'b00000_000000_00000;
		4138: oled_colour = 16'b00000_000000_00000;
		4139: oled_colour = 16'b00000_000000_00000;
		4140: oled_colour = 16'b00000_000000_00000;
		4141: oled_colour = 16'b00000_000000_00000;
		4142: oled_colour = 16'b00000_000000_00000;
		4143: oled_colour = 16'b00000_000000_00000;
		4144: oled_colour = 16'b00000_000000_00000;
		4145: oled_colour = 16'b00000_000000_00000;
		4146: oled_colour = 16'b00000_000000_00000;
		4147: oled_colour = 16'b00000_000000_00000;
		4148: oled_colour = 16'b00000_000000_00000;
		4149: oled_colour = 16'b00000_000000_00000;
		4150: oled_colour = 16'b00000_000000_00000;
		4151: oled_colour = 16'b00000_000000_00000;
		4152: oled_colour = 16'b00000_000000_00000;
		4153: oled_colour = 16'b00000_000000_00000;
		4154: oled_colour = 16'b00000_000000_00000;
		4155: oled_colour = 16'b00000_000000_00000;
		4156: oled_colour = 16'b00000_000000_00000;
		4157: oled_colour = 16'b00000_000000_00000;
		4158: oled_colour = 16'b00000_000000_00000;
		4159: oled_colour = 16'b00000_000000_00000;
		4160: oled_colour = 16'b00000_000000_00000;
		4161: oled_colour = 16'b00000_000000_00000;
		4162: oled_colour = 16'b00000_000000_00000;
		4163: oled_colour = 16'b00000_000000_00000;
		4164: oled_colour = 16'b00000_000000_00000;
		4165: oled_colour = 16'b00000_000000_00000;
		4166: oled_colour = 16'b00000_000000_00000;
		4167: oled_colour = 16'b00000_000000_00000;
		4168: oled_colour = 16'b00000_000000_00000;
		4169: oled_colour = 16'b00000_000000_00000;
		4170: oled_colour = 16'b00000_000000_00000;
		4171: oled_colour = 16'b11111_111111_11111; 
		4172: oled_colour = 16'b00000_000000_00000;
		4173: oled_colour = 16'b11011_110001_10111; 
		4174: oled_colour = 16'b11001_100010_01100; 
		4175: oled_colour = 16'b11001_100100_01110; 
		4176: oled_colour = 16'b11011_101100_10100; 
		4177: oled_colour = 16'b11100_101111_10100; 
		4178: oled_colour = 16'b11111_111001_11100; 
		4179: oled_colour = 16'b00000_000000_00000;
		4180: oled_colour = 16'b11111_111111_11111; 
		4181: oled_colour = 16'b00000_000000_00000;
		4182: oled_colour = 16'b00000_000000_00000;
		4183: oled_colour = 16'b00000_000000_00000;
		4184: oled_colour = 16'b00000_000000_00000;
		4185: oled_colour = 16'b00000_000000_00000;
		4186: oled_colour = 16'b00000_000000_00000;
		4187: oled_colour = 16'b00000_000000_00000;
		4188: oled_colour = 16'b00000_000000_00000;
		4189: oled_colour = 16'b00000_000000_00000;
		4190: oled_colour = 16'b00000_000000_00000;
		4191: oled_colour = 16'b00000_000000_00000;
		4192: oled_colour = 16'b00000_000000_00000;
		4193: oled_colour = 16'b00000_000000_00000;
		4194: oled_colour = 16'b00000_000000_00000;
		4195: oled_colour = 16'b00000_000000_00000;
		4196: oled_colour = 16'b00000_000000_00000;
		4197: oled_colour = 16'b00000_000000_00000;
		4198: oled_colour = 16'b00000_000000_00000;
		4199: oled_colour = 16'b00000_000000_00000;
		4200: oled_colour = 16'b00000_000000_00000;
		4201: oled_colour = 16'b00000_000000_00000;
		4202: oled_colour = 16'b00000_000000_00000;
		4203: oled_colour = 16'b00000_000000_00000;
		4204: oled_colour = 16'b00000_000000_00000;
		4205: oled_colour = 16'b00000_000000_00000;
		4206: oled_colour = 16'b00000_000000_00000;
		4207: oled_colour = 16'b00000_000000_00000;
		4208: oled_colour = 16'b00000_000000_00000;
		4209: oled_colour = 16'b00000_000000_00000;
		4210: oled_colour = 16'b00000_000000_00000;
		4211: oled_colour = 16'b00000_000000_00000;
		4212: oled_colour = 16'b00000_000000_00000;
		4213: oled_colour = 16'b00000_000000_00000;
		4214: oled_colour = 16'b00000_000000_00000;
		4215: oled_colour = 16'b00000_000000_00000;
		4216: oled_colour = 16'b00000_000000_00000;
		4217: oled_colour = 16'b00000_000000_00000;
		4218: oled_colour = 16'b00000_000000_00000;
		4219: oled_colour = 16'b00000_000000_00000;
		4220: oled_colour = 16'b00000_000000_00000;
		4221: oled_colour = 16'b00000_000000_00000;
		4222: oled_colour = 16'b00000_000000_00000;
		4223: oled_colour = 16'b00000_000000_00000;
		4224: oled_colour = 16'b00000_000000_00000;
		4225: oled_colour = 16'b00000_000000_00000;
		4226: oled_colour = 16'b00000_000000_00000;
		4227: oled_colour = 16'b00000_000000_00000;
		4228: oled_colour = 16'b00000_000000_00000;
		4229: oled_colour = 16'b00000_000000_00000;
		4230: oled_colour = 16'b00000_000000_00000;
		4231: oled_colour = 16'b00000_000000_00000;
		4232: oled_colour = 16'b00000_000000_00000;
		4233: oled_colour = 16'b00000_000000_00000;
		4234: oled_colour = 16'b00000_000000_00000;
		4235: oled_colour = 16'b00000_000000_00000;
		4236: oled_colour = 16'b00000_000000_00000;
		4237: oled_colour = 16'b00000_000000_00000;
		4238: oled_colour = 16'b00000_000000_00000;
		4239: oled_colour = 16'b00000_000000_00000;
		4240: oled_colour = 16'b00000_000000_00000;
		4241: oled_colour = 16'b00000_000000_00000;
		4242: oled_colour = 16'b00000_000000_00000;
		4243: oled_colour = 16'b00000_000000_00000;
		4244: oled_colour = 16'b00000_000000_00000;
		4245: oled_colour = 16'b00000_000000_00000;
		4246: oled_colour = 16'b00000_000000_00000;
		4247: oled_colour = 16'b00000_000000_00000;
		4248: oled_colour = 16'b00000_000000_00000;
		4249: oled_colour = 16'b00000_000000_00000;
		4250: oled_colour = 16'b00000_000000_00000;
		4251: oled_colour = 16'b00000_000000_00000;
		4252: oled_colour = 16'b00000_000000_00000;
		4253: oled_colour = 16'b00000_000000_00000;
		4254: oled_colour = 16'b00000_000000_00000;
		4255: oled_colour = 16'b00000_000000_00000;
		4256: oled_colour = 16'b00000_000000_00000;
		4257: oled_colour = 16'b00000_000000_00000;
		4258: oled_colour = 16'b00000_000000_00000;
		4259: oled_colour = 16'b00000_000000_00000;
		4260: oled_colour = 16'b00000_000000_00000;
		4261: oled_colour = 16'b00000_000000_00000;
		4262: oled_colour = 16'b00000_000000_00000;
		4263: oled_colour = 16'b00000_000000_00000;
		4264: oled_colour = 16'b00000_000000_00000;
		4265: oled_colour = 16'b00000_000000_00000;
		4266: oled_colour = 16'b00000_000000_00000;
		4267: oled_colour = 16'b00000_000000_00000;
		4268: oled_colour = 16'b00000_000000_00000;
		4269: oled_colour = 16'b11111_111111_11111; 
		4270: oled_colour = 16'b11101_110110_11010; 
		4271: oled_colour = 16'b11111_111010_11100; 
		4272: oled_colour = 16'b00000_000000_00000;
		4273: oled_colour = 16'b11111_111111_11111; 
		4274: oled_colour = 16'b00000_000000_00000;
		4275: oled_colour = 16'b00000_000000_00000;
		4276: oled_colour = 16'b00000_000000_00000;
		4277: oled_colour = 16'b00000_000000_00000;
		4278: oled_colour = 16'b00000_000000_00000;
		4279: oled_colour = 16'b00000_000000_00000;
		4280: oled_colour = 16'b00000_000000_00000;
		4281: oled_colour = 16'b00000_000000_00000;
		4282: oled_colour = 16'b00000_000000_00000;
		4283: oled_colour = 16'b00000_000000_00000;
		4284: oled_colour = 16'b00000_000000_00000;
		4285: oled_colour = 16'b00000_000000_00000;
		4286: oled_colour = 16'b00000_000000_00000;
		4287: oled_colour = 16'b00000_000000_00000;
		4288: oled_colour = 16'b00000_000000_00000;
		4289: oled_colour = 16'b00000_000000_00000;
		4290: oled_colour = 16'b00000_000000_00000;
		4291: oled_colour = 16'b00000_000000_00000;
		4292: oled_colour = 16'b00000_000000_00000;
		4293: oled_colour = 16'b00000_000000_00000;
		4294: oled_colour = 16'b00000_000000_00000;
		4295: oled_colour = 16'b00000_000000_00000;
		4296: oled_colour = 16'b00000_000000_00000;
		4297: oled_colour = 16'b00000_000000_00000;
		4298: oled_colour = 16'b00000_000000_00000;
		4299: oled_colour = 16'b00000_000000_00000;
		4300: oled_colour = 16'b00000_000000_00000;
		4301: oled_colour = 16'b00000_000000_00000;
		4302: oled_colour = 16'b00000_000000_00000;
		4303: oled_colour = 16'b00000_000000_00000;
		4304: oled_colour = 16'b00000_000000_00000;
		4305: oled_colour = 16'b00000_000000_00000;
		4306: oled_colour = 16'b00000_000000_00000;
		4307: oled_colour = 16'b00000_000000_00000;
		4308: oled_colour = 16'b00000_000000_00000;
		4309: oled_colour = 16'b00000_000000_00000;
		4310: oled_colour = 16'b00000_000000_00000;
		4311: oled_colour = 16'b00000_000000_00000;
		4312: oled_colour = 16'b00000_000000_00000;
		4313: oled_colour = 16'b00000_000000_00000;
		4314: oled_colour = 16'b00000_000000_00000;
		4315: oled_colour = 16'b00000_000000_00000;
		4316: oled_colour = 16'b00000_000000_00000;
		4317: oled_colour = 16'b00000_000000_00000;
		4318: oled_colour = 16'b00000_000000_00000;
		4319: oled_colour = 16'b00000_000000_00000;
		4320: oled_colour = 16'b00000_000000_00000;
		4321: oled_colour = 16'b00000_000000_00000;
		4322: oled_colour = 16'b00000_000000_00000;
		4323: oled_colour = 16'b00000_000000_00000;
		4324: oled_colour = 16'b00000_000000_00000;
		4325: oled_colour = 16'b00000_000000_00000;
		4326: oled_colour = 16'b00000_000000_00000;
		4327: oled_colour = 16'b00000_000000_00000;
		4328: oled_colour = 16'b00000_000000_00000;
		4329: oled_colour = 16'b00000_000000_00000;
		4330: oled_colour = 16'b00000_000000_00000;
		4331: oled_colour = 16'b00000_000000_00000;
		4332: oled_colour = 16'b00000_000000_00000;
		4333: oled_colour = 16'b00000_000000_00000;
		4334: oled_colour = 16'b00000_000000_00000;
		4335: oled_colour = 16'b00000_000000_00000;
		4336: oled_colour = 16'b00000_000000_00000;
		4337: oled_colour = 16'b00000_000000_00000;
		4338: oled_colour = 16'b00000_000000_00000;
		4339: oled_colour = 16'b00000_000000_00000;
		4340: oled_colour = 16'b00000_000000_00000;
		4341: oled_colour = 16'b00000_000000_00000;
		4342: oled_colour = 16'b00000_000000_00000;
		4343: oled_colour = 16'b00000_000000_00000;
		4344: oled_colour = 16'b00000_000000_00000;
		4345: oled_colour = 16'b00000_000000_00000;
		4346: oled_colour = 16'b00000_000000_00000;
		4347: oled_colour = 16'b00000_000000_00000;
		4348: oled_colour = 16'b00000_000000_00000;
		4349: oled_colour = 16'b00000_000000_00000;
		4350: oled_colour = 16'b00000_000000_00000;
		4351: oled_colour = 16'b00000_000000_00000;
		4352: oled_colour = 16'b00000_000000_00000;
		4353: oled_colour = 16'b00000_000000_00000;
		4354: oled_colour = 16'b00000_000000_00000;
		4355: oled_colour = 16'b00000_000000_00000;
		4356: oled_colour = 16'b00000_000000_00000;
		4357: oled_colour = 16'b00000_000000_00000;
		4358: oled_colour = 16'b00000_000000_00000;
		4359: oled_colour = 16'b00000_000000_00000;
		4360: oled_colour = 16'b00000_000000_00000;
		4361: oled_colour = 16'b00000_000000_00000;
		4362: oled_colour = 16'b00000_000000_00000;
		4363: oled_colour = 16'b00000_000000_00000;
		4364: oled_colour = 16'b00000_000000_00000;
		4365: oled_colour = 16'b00000_000000_00000;
		4366: oled_colour = 16'b00000_000000_00000;
		4367: oled_colour = 16'b00000_000000_00000;
		4368: oled_colour = 16'b00000_000000_00000;
		4369: oled_colour = 16'b00000_000000_00000;
		4370: oled_colour = 16'b11111_111111_11111; 
		4371: oled_colour = 16'b00000_000000_00000;
		4372: oled_colour = 16'b00000_000000_00000;
		4373: oled_colour = 16'b00000_000000_00000;
		4374: oled_colour = 16'b00000_000000_00000;
		4375: oled_colour = 16'b00000_000000_00000;
		4376: oled_colour = 16'b00000_000000_00000;
		4377: oled_colour = 16'b00000_000000_00000;
		4378: oled_colour = 16'b00000_000000_00000;
		4379: oled_colour = 16'b00000_000000_00000;
		4380: oled_colour = 16'b00000_000000_00000;
		4381: oled_colour = 16'b00000_000000_00000;
		4382: oled_colour = 16'b00000_000000_00000;
		4383: oled_colour = 16'b00000_000000_00000;
		4384: oled_colour = 16'b00000_000000_00000;
		4385: oled_colour = 16'b00000_000000_00000;
		4386: oled_colour = 16'b00000_000000_00000;
		4387: oled_colour = 16'b00000_000000_00000;
		4388: oled_colour = 16'b00000_000000_00000;
		4389: oled_colour = 16'b00000_000000_00000;
		4390: oled_colour = 16'b00000_000000_00000;
		4391: oled_colour = 16'b00000_000000_00000;
		4392: oled_colour = 16'b00000_000000_00000;
		4393: oled_colour = 16'b00000_000000_00000;
		4394: oled_colour = 16'b00000_000000_00000;
		4395: oled_colour = 16'b00000_000000_00000;
		4396: oled_colour = 16'b00000_000000_00000;
		4397: oled_colour = 16'b00000_000000_00000;
		4398: oled_colour = 16'b00000_000000_00000;
		4399: oled_colour = 16'b00000_000000_00000;
		4400: oled_colour = 16'b00000_000000_00000;
		4401: oled_colour = 16'b00000_000000_00000;
		4402: oled_colour = 16'b00000_000000_00000;
		4403: oled_colour = 16'b00000_000000_00000;
		4404: oled_colour = 16'b00000_000000_00000;
		4405: oled_colour = 16'b00000_000000_00000;
		4406: oled_colour = 16'b00000_000000_00000;
		4407: oled_colour = 16'b00000_000000_00000;
		4408: oled_colour = 16'b00000_000000_00000;
		4409: oled_colour = 16'b00000_000000_00000;
		4410: oled_colour = 16'b00000_000000_00000;
		4411: oled_colour = 16'b00000_000000_00000;
		4412: oled_colour = 16'b00000_000000_00000;
		4413: oled_colour = 16'b00000_000000_00000;
		4414: oled_colour = 16'b00000_000000_00000;
		4415: oled_colour = 16'b00000_000000_00000;
		4416: oled_colour = 16'b00000_000000_00000;
		4417: oled_colour = 16'b00000_000000_00000;
		4418: oled_colour = 16'b00000_000000_00000;
		4419: oled_colour = 16'b00000_000000_00000;
		4420: oled_colour = 16'b00000_000000_00000;
		4421: oled_colour = 16'b00000_000000_00000;
		4422: oled_colour = 16'b00000_000000_00000;
		4423: oled_colour = 16'b00000_000000_00000;
		4424: oled_colour = 16'b00000_000000_00000;
		4425: oled_colour = 16'b00000_000000_00000;
		4426: oled_colour = 16'b00000_000000_00000;
		4427: oled_colour = 16'b00000_000000_00000;
		4428: oled_colour = 16'b00000_000000_00000;
		4429: oled_colour = 16'b00000_000000_00000;
		4430: oled_colour = 16'b00000_000000_00000;
		4431: oled_colour = 16'b00000_000000_00000;
		4432: oled_colour = 16'b00000_000000_00000;
		4433: oled_colour = 16'b00000_000000_00000;
		4434: oled_colour = 16'b00000_000000_00000;
		4435: oled_colour = 16'b00000_000000_00000;
		4436: oled_colour = 16'b00000_000000_00000;
		4437: oled_colour = 16'b00000_000000_00000;
		4438: oled_colour = 16'b00000_000000_00000;
		4439: oled_colour = 16'b00000_000000_00000;
		4440: oled_colour = 16'b00000_000000_00000;
		4441: oled_colour = 16'b00000_000000_00000;
		4442: oled_colour = 16'b00000_000000_00000;
		4443: oled_colour = 16'b00000_000000_00000;
		4444: oled_colour = 16'b00000_000000_00000;
		4445: oled_colour = 16'b00000_000000_00000;
		4446: oled_colour = 16'b00000_000000_00000;
		4447: oled_colour = 16'b00000_000000_00000;
		4448: oled_colour = 16'b00000_000000_00000;
		4449: oled_colour = 16'b00000_000000_00000;
		4450: oled_colour = 16'b00000_000000_00000;
		4451: oled_colour = 16'b00000_000000_00000;
		4452: oled_colour = 16'b00000_000000_00000;
		4453: oled_colour = 16'b00000_000000_00000;
		4454: oled_colour = 16'b00000_000000_00000;
		4455: oled_colour = 16'b00000_000000_00000;
		4456: oled_colour = 16'b00000_000000_00000;
		4457: oled_colour = 16'b00000_000000_00000;
		4458: oled_colour = 16'b00000_000000_00000;
		4459: oled_colour = 16'b00000_000000_00000;
		4460: oled_colour = 16'b00000_000000_00000;
		4461: oled_colour = 16'b00000_000000_00000;
		4462: oled_colour = 16'b11111_111111_11111; 
		4463: oled_colour = 16'b11111_111111_11111; 
		4464: oled_colour = 16'b00000_000000_00000;
		4465: oled_colour = 16'b00000_000000_00000;
		4466: oled_colour = 16'b00000_000000_00000;
		4467: oled_colour = 16'b00000_000000_00000;
		4468: oled_colour = 16'b00000_000000_00000;
		4469: oled_colour = 16'b00000_000000_00000;
		4470: oled_colour = 16'b00000_000000_00000;
		4471: oled_colour = 16'b00000_000000_00000;
		4472: oled_colour = 16'b00000_000000_00000;
		4473: oled_colour = 16'b00000_000000_00000;
		4474: oled_colour = 16'b00000_000000_00000;
		4475: oled_colour = 16'b00000_000000_00000;
		4476: oled_colour = 16'b00000_000000_00000;
		4477: oled_colour = 16'b00000_000000_00000;
		4478: oled_colour = 16'b00000_000000_00000;
		4479: oled_colour = 16'b00000_000000_00000;
		4480: oled_colour = 16'b00000_000000_00000;
		4481: oled_colour = 16'b00000_000000_00000;
		4482: oled_colour = 16'b00000_000000_00000;
		4483: oled_colour = 16'b00000_000000_00000;
		4484: oled_colour = 16'b00000_000000_00000;
		4485: oled_colour = 16'b00000_000000_00000;
		4486: oled_colour = 16'b00000_000000_00000;
		4487: oled_colour = 16'b00000_000000_00000;
		4488: oled_colour = 16'b00000_000000_00000;
		4489: oled_colour = 16'b00000_000000_00000;
		4490: oled_colour = 16'b00000_000000_00000;
		4491: oled_colour = 16'b00000_000000_00000;
		4492: oled_colour = 16'b00000_000000_00000;
		4493: oled_colour = 16'b00000_000000_00000;
		4494: oled_colour = 16'b00000_000000_00000;
		4495: oled_colour = 16'b00000_000000_00000;
		4496: oled_colour = 16'b00000_000000_00000;
		4497: oled_colour = 16'b00000_000000_00000;
		4498: oled_colour = 16'b00000_000000_00000;
		4499: oled_colour = 16'b00000_000000_00000;
		4500: oled_colour = 16'b00000_000000_00000;
		4501: oled_colour = 16'b00000_000000_00000;
		4502: oled_colour = 16'b00000_000000_00000;
		4503: oled_colour = 16'b00000_000000_00000;
		4504: oled_colour = 16'b00000_000000_00000;
		4505: oled_colour = 16'b00000_000000_00000;
		4506: oled_colour = 16'b00000_000000_00000;
		4507: oled_colour = 16'b00000_000000_00000;
		4508: oled_colour = 16'b00000_000000_00000;
		4509: oled_colour = 16'b00000_000000_00000;
		4510: oled_colour = 16'b00000_000000_00000;
		4511: oled_colour = 16'b00000_000000_00000;
		4512: oled_colour = 16'b00000_000000_00000;
		4513: oled_colour = 16'b00000_000000_00000;
		4514: oled_colour = 16'b00000_000000_00000;
		4515: oled_colour = 16'b00000_000000_00000;
		4516: oled_colour = 16'b00000_000000_00000;
		4517: oled_colour = 16'b00000_000000_00000;
		4518: oled_colour = 16'b00000_000000_00000;
		4519: oled_colour = 16'b00000_000000_00000;
		4520: oled_colour = 16'b00000_000000_00000;
		4521: oled_colour = 16'b00000_000000_00000;
		4522: oled_colour = 16'b00000_000000_00000;
		4523: oled_colour = 16'b00000_000000_00000;
		4524: oled_colour = 16'b00000_000000_00000;
		4525: oled_colour = 16'b00000_000000_00000;
		4526: oled_colour = 16'b00000_000000_00000;
		4527: oled_colour = 16'b00000_000000_00000;
		4528: oled_colour = 16'b00000_000000_00000;
		4529: oled_colour = 16'b00000_000000_00000;
		4530: oled_colour = 16'b00000_000000_00000;
		4531: oled_colour = 16'b00000_000000_00000;
		4532: oled_colour = 16'b00000_000000_00000;
		4533: oled_colour = 16'b00000_000000_00000;
		4534: oled_colour = 16'b00000_000000_00000;
		4535: oled_colour = 16'b00000_000000_00000;
		4536: oled_colour = 16'b00000_000000_00000;
		4537: oled_colour = 16'b00000_000000_00000;
		4538: oled_colour = 16'b00000_000000_00000;
		4539: oled_colour = 16'b00000_000000_00000;
		4540: oled_colour = 16'b00000_000000_00000;
		4541: oled_colour = 16'b00000_000000_00000;
		4542: oled_colour = 16'b00000_000000_00000;
		4543: oled_colour = 16'b00000_000000_00000;
		4544: oled_colour = 16'b00000_000000_00000;
		4545: oled_colour = 16'b00000_000000_00000;
		4546: oled_colour = 16'b00000_000000_00000;
		4547: oled_colour = 16'b00000_000000_00000;
		4548: oled_colour = 16'b00000_000000_00000;
		4549: oled_colour = 16'b00000_000000_00000;
		4550: oled_colour = 16'b00000_000000_00000;
		4551: oled_colour = 16'b00000_000000_00000;
		4552: oled_colour = 16'b00000_000000_00000;
		4553: oled_colour = 16'b00000_000000_00000;
		4554: oled_colour = 16'b00000_000000_00000;
		4555: oled_colour = 16'b00000_000000_00000;
		4556: oled_colour = 16'b00000_000000_00000;
		4557: oled_colour = 16'b00000_000000_00000;
		4558: oled_colour = 16'b00000_000000_00000;
		4559: oled_colour = 16'b00000_000000_00000;
		4560: oled_colour = 16'b00000_000000_00000;
		4561: oled_colour = 16'b00000_000000_00000;
		4562: oled_colour = 16'b00000_000000_00000;
		4563: oled_colour = 16'b00000_000000_00000;
		4564: oled_colour = 16'b00000_000000_00000;
		4565: oled_colour = 16'b00000_000000_00000;
		4566: oled_colour = 16'b00000_000000_00000;
		4567: oled_colour = 16'b00000_000000_00000;
		4568: oled_colour = 16'b00000_000000_00000;
		4569: oled_colour = 16'b00000_000000_00000;
		4570: oled_colour = 16'b00000_000000_00000;
		4571: oled_colour = 16'b00000_000000_00000;
		4572: oled_colour = 16'b00000_000000_00000;
		4573: oled_colour = 16'b00000_000000_00000;
		4574: oled_colour = 16'b00000_000000_00000;
		4575: oled_colour = 16'b00000_000000_00000;
		4576: oled_colour = 16'b00000_000000_00000;
		4577: oled_colour = 16'b00000_000000_00000;
		4578: oled_colour = 16'b00000_000000_00000;
		4579: oled_colour = 16'b00000_000000_00000;
		4580: oled_colour = 16'b00000_000000_00000;
		4581: oled_colour = 16'b00000_000000_00000;
		4582: oled_colour = 16'b00000_000000_00000;
		4583: oled_colour = 16'b00000_000000_00000;
		4584: oled_colour = 16'b00000_000000_00000;
		4585: oled_colour = 16'b00000_000000_00000;
		4586: oled_colour = 16'b00000_000000_00000;
		4587: oled_colour = 16'b00000_000000_00000;
		4588: oled_colour = 16'b00000_000000_00000;
		4589: oled_colour = 16'b00000_000000_00000;
		4590: oled_colour = 16'b00000_000000_00000;
		4591: oled_colour = 16'b00000_000000_00000;
		4592: oled_colour = 16'b00000_000000_00000;
		4593: oled_colour = 16'b00000_000000_00000;
		4594: oled_colour = 16'b00000_000000_00000;
		4595: oled_colour = 16'b00000_000000_00000;
		4596: oled_colour = 16'b00000_000000_00000;
		4597: oled_colour = 16'b00000_000000_00000;
		4598: oled_colour = 16'b00000_000000_00000;
		4599: oled_colour = 16'b00000_000000_00000;
		4600: oled_colour = 16'b00000_000000_00000;
		4601: oled_colour = 16'b00000_000000_00000;
		4602: oled_colour = 16'b00000_000000_00000;
		4603: oled_colour = 16'b00000_000000_00000;
		4604: oled_colour = 16'b00000_000000_00000;
		4605: oled_colour = 16'b00000_000000_00000;
		4606: oled_colour = 16'b00000_000000_00000;
		4607: oled_colour = 16'b00000_000000_00000;
		4608: oled_colour = 16'b00000_000000_00000;
		4609: oled_colour = 16'b00000_000000_00000;
		4610: oled_colour = 16'b00000_000000_00000;
		4611: oled_colour = 16'b00000_000000_00000;
		4612: oled_colour = 16'b00000_000000_00000;
		4613: oled_colour = 16'b00000_000000_00000;
		4614: oled_colour = 16'b00000_000000_00000;
		4615: oled_colour = 16'b00000_000000_00000;
		4616: oled_colour = 16'b00000_000000_00000;
		4617: oled_colour = 16'b00000_000000_00000;
		4618: oled_colour = 16'b00000_000000_00000;
		4619: oled_colour = 16'b00000_000000_00000;
		4620: oled_colour = 16'b00000_000000_00000;
		4621: oled_colour = 16'b00000_000000_00000;
		4622: oled_colour = 16'b00000_000000_00000;
		4623: oled_colour = 16'b00000_000000_00000;
		4624: oled_colour = 16'b00000_000000_00000;
		4625: oled_colour = 16'b00000_000000_00000;
		4626: oled_colour = 16'b00000_000000_00000;
		4627: oled_colour = 16'b00000_000000_00000;
		4628: oled_colour = 16'b00000_000000_00000;
		4629: oled_colour = 16'b00000_000000_00000;
		4630: oled_colour = 16'b00000_000000_00000;
		4631: oled_colour = 16'b00000_000000_00000;
		4632: oled_colour = 16'b00000_000000_00000;
		4633: oled_colour = 16'b00000_000000_00000;
		4634: oled_colour = 16'b00000_000000_00000;
		4635: oled_colour = 16'b00000_000000_00000;
		4636: oled_colour = 16'b00000_000000_00000;
		4637: oled_colour = 16'b00000_000000_00000;
		4638: oled_colour = 16'b00000_000000_00000;
		4639: oled_colour = 16'b00000_000000_00000;
		4640: oled_colour = 16'b00000_000000_00000;
		4641: oled_colour = 16'b00000_000000_00000;
		4642: oled_colour = 16'b00000_000000_00000;
		4643: oled_colour = 16'b00000_000000_00000;
		4644: oled_colour = 16'b00000_000000_00000;
		4645: oled_colour = 16'b00000_000000_00000;
		4646: oled_colour = 16'b00000_000000_00000;
		4647: oled_colour = 16'b00000_000000_00000;
		4648: oled_colour = 16'b00000_000000_00000;
		4649: oled_colour = 16'b00000_000000_00000;
		4650: oled_colour = 16'b00000_000000_00000;
		4651: oled_colour = 16'b00000_000000_00000;
		4652: oled_colour = 16'b00000_000000_00000;
		4653: oled_colour = 16'b00000_000000_00000;
		4654: oled_colour = 16'b00000_000000_00000;
		4655: oled_colour = 16'b00000_000000_00000;
		4656: oled_colour = 16'b00000_000000_00000;
		4657: oled_colour = 16'b00000_000000_00000;
		4658: oled_colour = 16'b00000_000000_00000;
		4659: oled_colour = 16'b00000_000000_00000;
		4660: oled_colour = 16'b00000_000000_00000;
		4661: oled_colour = 16'b00000_000000_00000;
		4662: oled_colour = 16'b00000_000000_00000;
		4663: oled_colour = 16'b00000_000000_00000;
		4664: oled_colour = 16'b00000_000000_00000;
		4665: oled_colour = 16'b00000_000000_00000;
		4666: oled_colour = 16'b00000_000000_00000;
		4667: oled_colour = 16'b00000_000000_00000;
		4668: oled_colour = 16'b00000_000000_00000;
		4669: oled_colour = 16'b00000_000000_00000;
		4670: oled_colour = 16'b00000_000000_00000;
		4671: oled_colour = 16'b00000_000000_00000;
		4672: oled_colour = 16'b00000_000000_00000;
		4673: oled_colour = 16'b00000_000000_00000;
		4674: oled_colour = 16'b00000_000000_00000;
		4675: oled_colour = 16'b00000_000000_00000;
		4676: oled_colour = 16'b00000_000000_00000;
		4677: oled_colour = 16'b00000_000000_00000;
		4678: oled_colour = 16'b00000_000000_00000;
		4679: oled_colour = 16'b00000_000000_00000;
		4680: oled_colour = 16'b00000_000000_00000;
		4681: oled_colour = 16'b00000_000000_00000;
		4682: oled_colour = 16'b00000_000000_00000;
		4683: oled_colour = 16'b00000_000000_00000;
		4684: oled_colour = 16'b00000_000000_00000;
		4685: oled_colour = 16'b00000_000000_00000;
		4686: oled_colour = 16'b00000_000000_00000;
		4687: oled_colour = 16'b00000_000000_00000;
		4688: oled_colour = 16'b00000_000000_00000;
		4689: oled_colour = 16'b00000_000000_00000;
		4690: oled_colour = 16'b00000_000000_00000;
		4691: oled_colour = 16'b00000_000000_00000;
		4692: oled_colour = 16'b00000_000000_00000;
		4693: oled_colour = 16'b00000_000000_00000;
		4694: oled_colour = 16'b00000_000000_00000;
		4695: oled_colour = 16'b00000_000000_00000;
		4696: oled_colour = 16'b00000_000000_00000;
		4697: oled_colour = 16'b00000_000000_00000;
		4698: oled_colour = 16'b00000_000000_00000;
		4699: oled_colour = 16'b00000_000000_00000;
		4700: oled_colour = 16'b00000_000000_00000;
		4701: oled_colour = 16'b00000_000000_00000;
		4702: oled_colour = 16'b00000_000000_00000;
		4703: oled_colour = 16'b00000_000000_00000;
		4704: oled_colour = 16'b00000_000000_00000;
		4705: oled_colour = 16'b00000_000000_00000;
		4706: oled_colour = 16'b00000_000000_00000;
		4707: oled_colour = 16'b00000_000000_00000;
		4708: oled_colour = 16'b00000_000000_00000;
		4709: oled_colour = 16'b00000_000000_00000;
		4710: oled_colour = 16'b00000_000000_00000;
		4711: oled_colour = 16'b00000_000000_00000;
		4712: oled_colour = 16'b00000_000000_00000;
		4713: oled_colour = 16'b00000_000000_00000;
		4714: oled_colour = 16'b00000_000000_00000;
		4715: oled_colour = 16'b00000_000000_00000;
		4716: oled_colour = 16'b00000_000000_00000;
		4717: oled_colour = 16'b00000_000000_00000;
		4718: oled_colour = 16'b00000_000000_00000;
		4719: oled_colour = 16'b00000_000000_00000;
		4720: oled_colour = 16'b00000_000000_00000;
		4721: oled_colour = 16'b00000_000000_00000;
		4722: oled_colour = 16'b00000_000000_00000;
		4723: oled_colour = 16'b00000_000000_00000;
		4724: oled_colour = 16'b00000_000000_00000;
		4725: oled_colour = 16'b00000_000000_00000;
		4726: oled_colour = 16'b00000_000000_00000;
		4727: oled_colour = 16'b00000_000000_00000;
		4728: oled_colour = 16'b00000_000000_00000;
		4729: oled_colour = 16'b00000_000000_00000;
		4730: oled_colour = 16'b00000_000000_00000;
		4731: oled_colour = 16'b00000_000000_00000;
		4732: oled_colour = 16'b00000_000000_00000;
		4733: oled_colour = 16'b00000_000000_00000;
		4734: oled_colour = 16'b00000_000000_00000;
		4735: oled_colour = 16'b00000_000000_00000;
		4736: oled_colour = 16'b00000_000000_00000;
		4737: oled_colour = 16'b00000_000000_00000;
		4738: oled_colour = 16'b00000_000000_00000;
		4739: oled_colour = 16'b00000_000000_00000;
		4740: oled_colour = 16'b00000_000000_00000;
		4741: oled_colour = 16'b00000_000000_00000;
		4742: oled_colour = 16'b00000_000000_00000;
		4743: oled_colour = 16'b00000_000000_00000;
		4744: oled_colour = 16'b00000_000000_00000;
		4745: oled_colour = 16'b00000_000000_00000;
		4746: oled_colour = 16'b00000_000000_00000;
		4747: oled_colour = 16'b00000_000000_00000;
		4748: oled_colour = 16'b00000_000000_00000;
		4749: oled_colour = 16'b00000_000000_00000;
		4750: oled_colour = 16'b00000_000000_00000;
		4751: oled_colour = 16'b00000_000000_00000;
		4752: oled_colour = 16'b00000_000000_00000;
		4753: oled_colour = 16'b00000_000000_00000;
		4754: oled_colour = 16'b00000_000000_00000;
		4755: oled_colour = 16'b00000_000000_00000;
		4756: oled_colour = 16'b00000_000000_00000;
		4757: oled_colour = 16'b00000_000000_00000;
		4758: oled_colour = 16'b00000_000000_00000;
		4759: oled_colour = 16'b00000_000000_00000;
		4760: oled_colour = 16'b00000_000000_00000;
		4761: oled_colour = 16'b00000_000000_00000;
		4762: oled_colour = 16'b00000_000000_00000;
		4763: oled_colour = 16'b00000_000000_00000;
		4764: oled_colour = 16'b00000_000000_00000;
		4765: oled_colour = 16'b00000_000000_00000;
		4766: oled_colour = 16'b00000_000000_00000;
		4767: oled_colour = 16'b00000_000000_00000;
		4768: oled_colour = 16'b00000_000000_00000;
		4769: oled_colour = 16'b00000_000000_00000;
		4770: oled_colour = 16'b00000_000000_00000;
		4771: oled_colour = 16'b00000_000000_00000;
		4772: oled_colour = 16'b00000_000000_00000;
		4773: oled_colour = 16'b00000_000000_00000;
		4774: oled_colour = 16'b00000_000000_00000;
		4775: oled_colour = 16'b00000_000000_00000;
		4776: oled_colour = 16'b00000_000000_00000;
		4777: oled_colour = 16'b00000_000000_00000;
		4778: oled_colour = 16'b00000_000000_00000;
		4779: oled_colour = 16'b00000_000000_00000;
		4780: oled_colour = 16'b00000_000000_00000;
		4781: oled_colour = 16'b00000_000000_00000;
		4782: oled_colour = 16'b00000_000000_00000;
		4783: oled_colour = 16'b00000_000000_00000;
		4784: oled_colour = 16'b00000_000000_00000;
		4785: oled_colour = 16'b00000_000000_00000;
		4786: oled_colour = 16'b00000_000000_00000;
		4787: oled_colour = 16'b00000_000000_00000;
		4788: oled_colour = 16'b00000_000000_00000;
		4789: oled_colour = 16'b00000_000000_00000;
		4790: oled_colour = 16'b00000_000000_00000;
		4791: oled_colour = 16'b00000_000000_00000;
		4792: oled_colour = 16'b00000_000000_00000;
		4793: oled_colour = 16'b00000_000000_00000;
		4794: oled_colour = 16'b00000_000000_00000;
		4795: oled_colour = 16'b00000_000000_00000;
		4796: oled_colour = 16'b00000_000000_00000;
		4797: oled_colour = 16'b00000_000000_00000;
		4798: oled_colour = 16'b00000_000000_00000;
		4799: oled_colour = 16'b00000_000000_00000;
		4800: oled_colour = 16'b00000_000000_00000;
		4801: oled_colour = 16'b00000_000000_00000;
		4802: oled_colour = 16'b00000_000000_00000;
		4803: oled_colour = 16'b00000_000000_00000;
		4804: oled_colour = 16'b00000_000000_00000;
		4805: oled_colour = 16'b00000_000000_00000;
		4806: oled_colour = 16'b00000_000000_00000;
		4807: oled_colour = 16'b00000_000000_00000;
		4808: oled_colour = 16'b00000_000000_00000;
		4809: oled_colour = 16'b00000_000000_00000;
		4810: oled_colour = 16'b00000_000000_00000;
		4811: oled_colour = 16'b00000_000000_00000;
		4812: oled_colour = 16'b00000_000000_00000;
		4813: oled_colour = 16'b00000_000000_00000;
		4814: oled_colour = 16'b00000_000000_00000;
		4815: oled_colour = 16'b00000_000000_00000;
		4816: oled_colour = 16'b00000_000000_00000;
		4817: oled_colour = 16'b00000_000000_00000;
		4818: oled_colour = 16'b00000_000000_00000;
		4819: oled_colour = 16'b00000_000000_00000;
		4820: oled_colour = 16'b00000_000000_00000;
		4821: oled_colour = 16'b00000_000000_00000;
		4822: oled_colour = 16'b00000_000000_00000;
		4823: oled_colour = 16'b00000_000000_00000;
		4824: oled_colour = 16'b00000_000000_00000;
		4825: oled_colour = 16'b00000_000000_00000;
		4826: oled_colour = 16'b00000_000000_00000;
		4827: oled_colour = 16'b00000_000000_00000;
		4828: oled_colour = 16'b00000_000000_00000;
		4829: oled_colour = 16'b00000_000000_00000;
		4830: oled_colour = 16'b00000_000000_00000;
		4831: oled_colour = 16'b00000_000000_00000;
		4832: oled_colour = 16'b00000_000000_00000;
		4833: oled_colour = 16'b00000_000000_00000;
		4834: oled_colour = 16'b00000_000000_00000;
		4835: oled_colour = 16'b00000_000000_00000;
		4836: oled_colour = 16'b00000_000000_00000;
		4837: oled_colour = 16'b00000_000000_00000;
		4838: oled_colour = 16'b00000_000000_00000;
		4839: oled_colour = 16'b00000_000000_00000;
		4840: oled_colour = 16'b00000_000000_00000;
		4841: oled_colour = 16'b00000_000000_00000;
		4842: oled_colour = 16'b00000_000000_00000;
		4843: oled_colour = 16'b00000_000000_00000;
		4844: oled_colour = 16'b00000_000000_00000;
		4845: oled_colour = 16'b00000_000000_00000;
		4846: oled_colour = 16'b00000_000000_00000;
		4847: oled_colour = 16'b00000_000000_00000;
		4848: oled_colour = 16'b00000_000000_00000;
		4849: oled_colour = 16'b00000_000000_00000;
		4850: oled_colour = 16'b00000_000000_00000;
		4851: oled_colour = 16'b00000_000000_00000;
		4852: oled_colour = 16'b00000_000000_00000;
		4853: oled_colour = 16'b00000_000000_00000;
		4854: oled_colour = 16'b00000_000000_00000;
		4855: oled_colour = 16'b00000_000000_00000;
		4856: oled_colour = 16'b00000_000000_00000;
		4857: oled_colour = 16'b00000_000000_00000;
		4858: oled_colour = 16'b00000_000000_00000;
		4859: oled_colour = 16'b00000_000000_00000;
		4860: oled_colour = 16'b00000_000000_00000;
		4861: oled_colour = 16'b00000_000000_00000;
		4862: oled_colour = 16'b00000_000000_00000;
		4863: oled_colour = 16'b00000_000000_00000;
		4864: oled_colour = 16'b00000_000000_00000;
		4865: oled_colour = 16'b00000_000000_00000;
		4866: oled_colour = 16'b00000_000000_00000;
		4867: oled_colour = 16'b00000_000000_00000;
		4868: oled_colour = 16'b00000_000000_00000;
		4869: oled_colour = 16'b00000_000000_00000;
		4870: oled_colour = 16'b00000_000000_00000;
		4871: oled_colour = 16'b00000_000000_00000;
		4872: oled_colour = 16'b00000_000000_00000;
		4873: oled_colour = 16'b00000_000000_00000;
		4874: oled_colour = 16'b00000_000000_00000;
		4875: oled_colour = 16'b00000_000000_00000;
		4876: oled_colour = 16'b00000_000000_00000;
		4877: oled_colour = 16'b00000_000000_00000;
		4878: oled_colour = 16'b00000_000000_00000;
		4879: oled_colour = 16'b00000_000000_00000;
		4880: oled_colour = 16'b00000_000000_00000;
		4881: oled_colour = 16'b00000_000000_00000;
		4882: oled_colour = 16'b00000_000000_00000;
		4883: oled_colour = 16'b00000_000000_00000;
		4884: oled_colour = 16'b00000_000000_00000;
		4885: oled_colour = 16'b00000_000000_00000;
		4886: oled_colour = 16'b00000_000000_00000;
		4887: oled_colour = 16'b00000_000000_00000;
		4888: oled_colour = 16'b00000_000000_00000;
		4889: oled_colour = 16'b00000_000000_00000;
		4890: oled_colour = 16'b00000_000000_00000;
		4891: oled_colour = 16'b00000_000000_00000;
		4892: oled_colour = 16'b00000_000000_00000;
		4893: oled_colour = 16'b00000_000000_00000;
		4894: oled_colour = 16'b00000_000000_00000;
		4895: oled_colour = 16'b00000_000000_00000;
		4896: oled_colour = 16'b00000_000000_00000;
		4897: oled_colour = 16'b00000_000000_00000;
		4898: oled_colour = 16'b00000_000000_00000;
		4899: oled_colour = 16'b00000_000000_00000;
		4900: oled_colour = 16'b00000_000000_00000;
		4901: oled_colour = 16'b00000_000000_00000;
		4902: oled_colour = 16'b00000_000000_00000;
		4903: oled_colour = 16'b00000_000000_00000;
		4904: oled_colour = 16'b00000_000000_00000;
		4905: oled_colour = 16'b00000_000000_00000;
		4906: oled_colour = 16'b00000_000000_00000;
		4907: oled_colour = 16'b00000_000000_00000;
		4908: oled_colour = 16'b00000_000000_00000;
		4909: oled_colour = 16'b00000_000000_00000;
		4910: oled_colour = 16'b00000_000000_00000;
		4911: oled_colour = 16'b00000_000000_00000;
		4912: oled_colour = 16'b00000_000000_00000;
		4913: oled_colour = 16'b00000_000000_00000;
		4914: oled_colour = 16'b00000_000000_00000;
		4915: oled_colour = 16'b00000_000000_00000;
		4916: oled_colour = 16'b00000_000000_00000;
		4917: oled_colour = 16'b00000_000000_00000;
		4918: oled_colour = 16'b00000_000000_00000;
		4919: oled_colour = 16'b00000_000000_00000;
		4920: oled_colour = 16'b00000_000000_00000;
		4921: oled_colour = 16'b00000_000000_00000;
		4922: oled_colour = 16'b00000_000000_00000;
		4923: oled_colour = 16'b00000_000000_00000;
		4924: oled_colour = 16'b00000_000000_00000;
		4925: oled_colour = 16'b00000_000000_00000;
		4926: oled_colour = 16'b00000_000000_00000;
		4927: oled_colour = 16'b00000_000000_00000;
		4928: oled_colour = 16'b00000_000000_00000;
		4929: oled_colour = 16'b00000_000000_00000;
		4930: oled_colour = 16'b00000_000000_00000;
		4931: oled_colour = 16'b00000_000000_00000;
		4932: oled_colour = 16'b00000_000000_00000;
		4933: oled_colour = 16'b00000_000000_00000;
		4934: oled_colour = 16'b00000_000000_00000;
		4935: oled_colour = 16'b00000_000000_00000;
		4936: oled_colour = 16'b00000_000000_00000;
		4937: oled_colour = 16'b00000_000000_00000;
		4938: oled_colour = 16'b00000_000000_00000;
		4939: oled_colour = 16'b00000_000000_00000;
		4940: oled_colour = 16'b00000_000000_00000;
		4941: oled_colour = 16'b00000_000000_00000;
		4942: oled_colour = 16'b00000_000000_00000;
		4943: oled_colour = 16'b00000_000000_00000;
		4944: oled_colour = 16'b00000_000000_00000;
		4945: oled_colour = 16'b00000_000000_00000;
		4946: oled_colour = 16'b00000_000000_00000;
		4947: oled_colour = 16'b00000_000000_00000;
		4948: oled_colour = 16'b00000_000000_00000;
		4949: oled_colour = 16'b00000_000000_00000;
		4950: oled_colour = 16'b00000_000000_00000;
		4951: oled_colour = 16'b00000_000000_00000;
		4952: oled_colour = 16'b00000_000000_00000;
		4953: oled_colour = 16'b00000_000000_00000;
		4954: oled_colour = 16'b00000_000000_00000;
		4955: oled_colour = 16'b00000_000000_00000;
		4956: oled_colour = 16'b00000_000000_00000;
		4957: oled_colour = 16'b00000_000000_00000;
		4958: oled_colour = 16'b00000_000000_00000;
		4959: oled_colour = 16'b00000_000000_00000;
		4960: oled_colour = 16'b00000_000000_00000;
		4961: oled_colour = 16'b00000_000000_00000;
		4962: oled_colour = 16'b00000_000000_00000;
		4963: oled_colour = 16'b00000_000000_00000;
		4964: oled_colour = 16'b00000_000000_00000;
		4965: oled_colour = 16'b00000_000000_00000;
		4966: oled_colour = 16'b00000_000000_00000;
		4967: oled_colour = 16'b00000_000000_00000;
		4968: oled_colour = 16'b00000_000000_00000;
		4969: oled_colour = 16'b00000_000000_00000;
		4970: oled_colour = 16'b00000_000000_00000;
		4971: oled_colour = 16'b00000_000000_00000;
		4972: oled_colour = 16'b00000_000000_00000;
		4973: oled_colour = 16'b00000_000000_00000;
		4974: oled_colour = 16'b00000_000000_00000;
		4975: oled_colour = 16'b00000_000000_00000;
		4976: oled_colour = 16'b00000_000000_00000;
		4977: oled_colour = 16'b00000_000000_00000;
		4978: oled_colour = 16'b00000_000000_00000;
		4979: oled_colour = 16'b00000_000000_00000;
		4980: oled_colour = 16'b00000_000000_00000;
		4981: oled_colour = 16'b00000_000000_00000;
		4982: oled_colour = 16'b00000_000000_00000;
		4983: oled_colour = 16'b00000_000000_00000;
		4984: oled_colour = 16'b00000_000000_00000;
		4985: oled_colour = 16'b00000_000000_00000;
		4986: oled_colour = 16'b00000_000000_00000;
		4987: oled_colour = 16'b00000_000000_00000;
		4988: oled_colour = 16'b00000_000000_00000;
		4989: oled_colour = 16'b00000_000000_00000;
		4990: oled_colour = 16'b00000_000000_00000;
		4991: oled_colour = 16'b00000_000000_00000;
		4992: oled_colour = 16'b00000_000000_00000;
		4993: oled_colour = 16'b00000_000000_00000;
		4994: oled_colour = 16'b00000_000000_00000;
		4995: oled_colour = 16'b00000_000000_00000;
		4996: oled_colour = 16'b00000_000000_00000;
		4997: oled_colour = 16'b00000_000000_00000;
		4998: oled_colour = 16'b00000_000000_00000;
		4999: oled_colour = 16'b00000_000000_00000;
		5000: oled_colour = 16'b00000_000000_00000;
		5001: oled_colour = 16'b00000_000000_00000;
		5002: oled_colour = 16'b00000_000000_00000;
		5003: oled_colour = 16'b00000_000000_00000;
		5004: oled_colour = 16'b00000_000000_00000;
		5005: oled_colour = 16'b00000_000000_00000;
		5006: oled_colour = 16'b00000_000000_00000;
		5007: oled_colour = 16'b00000_000000_00000;
		5008: oled_colour = 16'b00000_000000_00000;
		5009: oled_colour = 16'b00000_000000_00000;
		5010: oled_colour = 16'b00000_000000_00000;
		5011: oled_colour = 16'b00000_000000_00000;
		5012: oled_colour = 16'b00000_000000_00000;
		5013: oled_colour = 16'b00000_000000_00000;
		5014: oled_colour = 16'b00000_000000_00000;
		5015: oled_colour = 16'b00000_000000_00000;
		5016: oled_colour = 16'b00000_000000_00000;
		5017: oled_colour = 16'b00000_000000_00000;
		5018: oled_colour = 16'b00000_000000_00000;
		5019: oled_colour = 16'b00000_000000_00000;
		5020: oled_colour = 16'b00000_000000_00000;
		5021: oled_colour = 16'b00000_000000_00000;
		5022: oled_colour = 16'b00000_000000_00000;
		5023: oled_colour = 16'b00000_000000_00000;
		5024: oled_colour = 16'b00000_000000_00000;
		5025: oled_colour = 16'b00000_000000_00000;
		5026: oled_colour = 16'b00000_000000_00000;
		5027: oled_colour = 16'b00000_000000_00000;
		5028: oled_colour = 16'b00000_000000_00000;
		5029: oled_colour = 16'b00000_000000_00000;
		5030: oled_colour = 16'b00000_000000_00000;
		5031: oled_colour = 16'b00000_000000_00000;
		5032: oled_colour = 16'b00000_000000_00000;
		5033: oled_colour = 16'b00000_000000_00000;
		5034: oled_colour = 16'b00000_000000_00000;
		5035: oled_colour = 16'b00000_000000_00000;
		5036: oled_colour = 16'b00000_000000_00000;
		5037: oled_colour = 16'b00000_000000_00000;
		5038: oled_colour = 16'b00000_000000_00000;
		5039: oled_colour = 16'b00000_000000_00000;
		5040: oled_colour = 16'b00000_000000_00000;
		5041: oled_colour = 16'b00000_000000_00000;
		5042: oled_colour = 16'b00000_000000_00000;
		5043: oled_colour = 16'b00000_000000_00000;
		5044: oled_colour = 16'b00000_000000_00000;
		5045: oled_colour = 16'b00000_000000_00000;
		5046: oled_colour = 16'b00000_000000_00000;
		5047: oled_colour = 16'b00000_000000_00000;
		5048: oled_colour = 16'b00000_000000_00000;
		5049: oled_colour = 16'b00000_000000_00000;
		5050: oled_colour = 16'b00000_000000_00000;
		5051: oled_colour = 16'b00000_000000_00000;
		5052: oled_colour = 16'b00000_000000_00000;
		5053: oled_colour = 16'b00000_000000_00000;
		5054: oled_colour = 16'b00000_000000_00000;
		5055: oled_colour = 16'b00000_000000_00000;
		5056: oled_colour = 16'b00000_000000_00000;
		5057: oled_colour = 16'b00000_000000_00000;
		5058: oled_colour = 16'b00000_000000_00000;
		5059: oled_colour = 16'b00000_000000_00000;
		5060: oled_colour = 16'b00000_000000_00000;
		5061: oled_colour = 16'b00000_000000_00000;
		5062: oled_colour = 16'b00000_000000_00000;
		5063: oled_colour = 16'b00000_000000_00000;
		5064: oled_colour = 16'b00000_000000_00000;
		5065: oled_colour = 16'b00000_000000_00000;
		5066: oled_colour = 16'b00000_000000_00000;
		5067: oled_colour = 16'b00000_000000_00000;
		5068: oled_colour = 16'b00000_000000_00000;
		5069: oled_colour = 16'b00000_000000_00000;
		5070: oled_colour = 16'b00000_000000_00000;
		5071: oled_colour = 16'b00000_000000_00000;
		5072: oled_colour = 16'b00000_000000_00000;
		5073: oled_colour = 16'b00000_000000_00000;
		5074: oled_colour = 16'b00000_000000_00000;
		5075: oled_colour = 16'b00000_000000_00000;
		5076: oled_colour = 16'b00000_000000_00000;
		5077: oled_colour = 16'b00000_000000_00000;
		5078: oled_colour = 16'b00000_000000_00000;
		5079: oled_colour = 16'b00000_000000_00000;
		5080: oled_colour = 16'b00000_000000_00000;
		5081: oled_colour = 16'b00000_000000_00000;
		5082: oled_colour = 16'b00000_000000_00000;
		5083: oled_colour = 16'b00000_000000_00000;
		5084: oled_colour = 16'b00000_000000_00000;
		5085: oled_colour = 16'b00000_000000_00000;
		5086: oled_colour = 16'b00000_000000_00000;
		5087: oled_colour = 16'b00000_000000_00000;
		5088: oled_colour = 16'b00000_000000_00000;
		5089: oled_colour = 16'b00000_000000_00000;
		5090: oled_colour = 16'b00000_000000_00000;
		5091: oled_colour = 16'b00000_000000_00000;
		5092: oled_colour = 16'b00000_000000_00000;
		5093: oled_colour = 16'b00000_000000_00000;
		5094: oled_colour = 16'b00000_000000_00000;
		5095: oled_colour = 16'b00000_000000_00000;
		5096: oled_colour = 16'b00000_000000_00000;
		5097: oled_colour = 16'b00000_000000_00000;
		5098: oled_colour = 16'b00000_000000_00000;
		5099: oled_colour = 16'b00000_000000_00000;
		5100: oled_colour = 16'b00000_000000_00000;
		5101: oled_colour = 16'b00000_000000_00000;
		5102: oled_colour = 16'b00000_000000_00000;
		5103: oled_colour = 16'b00000_000000_00000;
		5104: oled_colour = 16'b00000_000000_00000;
		5105: oled_colour = 16'b00000_000000_00000;
		5106: oled_colour = 16'b00000_000000_00000;
		5107: oled_colour = 16'b00000_000000_00000;
		5108: oled_colour = 16'b00000_000000_00000;
		5109: oled_colour = 16'b00000_000000_00000;
		5110: oled_colour = 16'b00000_000000_00000;
		5111: oled_colour = 16'b00000_000000_00000;
		5112: oled_colour = 16'b00000_000000_00000;
		5113: oled_colour = 16'b00000_000000_00000;
		5114: oled_colour = 16'b00000_000000_00000;
		5115: oled_colour = 16'b00000_000000_00000;
		5116: oled_colour = 16'b00000_000000_00000;
		5117: oled_colour = 16'b00000_000000_00000;
		5118: oled_colour = 16'b00000_000000_00000;
		5119: oled_colour = 16'b00000_000000_00000;
		5120: oled_colour = 16'b00000_000000_00000;
		5121: oled_colour = 16'b00000_000000_00000;
		5122: oled_colour = 16'b00000_000000_00000;
		5123: oled_colour = 16'b00000_000000_00000;
		5124: oled_colour = 16'b00000_000000_00000;
		5125: oled_colour = 16'b00000_000000_00000;
		5126: oled_colour = 16'b00000_000000_00000;
		5127: oled_colour = 16'b00000_000000_00000;
		5128: oled_colour = 16'b00000_000000_00000;
		5129: oled_colour = 16'b00000_000000_00000;
		5130: oled_colour = 16'b00000_000000_00000;
		5131: oled_colour = 16'b00000_000000_00000;
		5132: oled_colour = 16'b00000_000000_00000;
		5133: oled_colour = 16'b00000_000000_00000;
		5134: oled_colour = 16'b00000_000000_00000;
		5135: oled_colour = 16'b00000_000000_00000;
		5136: oled_colour = 16'b00000_000000_00000;
		5137: oled_colour = 16'b00000_000000_00000;
		5138: oled_colour = 16'b00000_000000_00000;
		5139: oled_colour = 16'b00000_000000_00000;
		5140: oled_colour = 16'b00000_000000_00000;
		5141: oled_colour = 16'b00000_000000_00000;
		5142: oled_colour = 16'b00000_000000_00000;
		5143: oled_colour = 16'b00000_000000_00000;
		5144: oled_colour = 16'b00000_000000_00000;
		5145: oled_colour = 16'b00000_000000_00000;
		5146: oled_colour = 16'b00000_000000_00000;
		5147: oled_colour = 16'b00000_000000_00000;
		5148: oled_colour = 16'b00000_000000_00000;
		5149: oled_colour = 16'b00000_000000_00000;
		5150: oled_colour = 16'b00000_000000_00000;
		5151: oled_colour = 16'b00000_000000_00000;
		5152: oled_colour = 16'b00000_000000_00000;
		5153: oled_colour = 16'b00000_000000_00000;
		5154: oled_colour = 16'b00000_000000_00000;
		5155: oled_colour = 16'b00000_000000_00000;
		5156: oled_colour = 16'b00000_000000_00000;
		5157: oled_colour = 16'b00000_000000_00000;
		5158: oled_colour = 16'b00000_000000_00000;
		5159: oled_colour = 16'b00000_000000_00000;
		5160: oled_colour = 16'b00000_000000_00000;
		5161: oled_colour = 16'b00000_000000_00000;
		5162: oled_colour = 16'b00000_000000_00000;
		5163: oled_colour = 16'b00000_000000_00000;
		5164: oled_colour = 16'b00000_000000_00000;
		5165: oled_colour = 16'b00000_000000_00000;
		5166: oled_colour = 16'b00000_000000_00000;
		5167: oled_colour = 16'b00000_000000_00000;
		5168: oled_colour = 16'b00000_000000_00000;
		5169: oled_colour = 16'b00000_000000_00000;
		5170: oled_colour = 16'b00000_000000_00000;
		5171: oled_colour = 16'b00000_000000_00000;
		5172: oled_colour = 16'b00000_000000_00000;
		5173: oled_colour = 16'b00000_000000_00000;
		5174: oled_colour = 16'b00000_000000_00000;
		5175: oled_colour = 16'b00000_000000_00000;
		5176: oled_colour = 16'b00000_000000_00000;
		5177: oled_colour = 16'b00000_000000_00000;
		5178: oled_colour = 16'b00000_000000_00000;
		5179: oled_colour = 16'b00000_000000_00000;
		5180: oled_colour = 16'b00000_000000_00000;
		5181: oled_colour = 16'b00000_000000_00000;
		5182: oled_colour = 16'b00000_000000_00000;
		5183: oled_colour = 16'b00000_000000_00000;
		5184: oled_colour = 16'b00000_000000_00000;
		5185: oled_colour = 16'b00000_000000_00000;
		5186: oled_colour = 16'b00000_000000_00000;
		5187: oled_colour = 16'b00000_000000_00000;
		5188: oled_colour = 16'b00000_000000_00000;
		5189: oled_colour = 16'b00000_000000_00000;
		5190: oled_colour = 16'b00000_000000_00000;
		5191: oled_colour = 16'b00000_000000_00000;
		5192: oled_colour = 16'b00000_000000_00000;
		5193: oled_colour = 16'b00000_000000_00000;
		5194: oled_colour = 16'b00000_000000_00000;
		5195: oled_colour = 16'b00000_000000_00000;
		5196: oled_colour = 16'b00000_000000_00000;
		5197: oled_colour = 16'b00000_000000_00000;
		5198: oled_colour = 16'b00000_000000_00000;
		5199: oled_colour = 16'b00000_000000_00000;
		5200: oled_colour = 16'b00000_000000_00000;
		5201: oled_colour = 16'b00000_000000_00000;
		5202: oled_colour = 16'b00000_000000_00000;
		5203: oled_colour = 16'b00000_000000_00000;
		5204: oled_colour = 16'b00000_000000_00000;
		5205: oled_colour = 16'b00000_000000_00000;
		5206: oled_colour = 16'b00000_000000_00000;
		5207: oled_colour = 16'b00000_000000_00000;
		5208: oled_colour = 16'b00000_000000_00000;
		5209: oled_colour = 16'b00000_000000_00000;
		5210: oled_colour = 16'b00000_000000_00000;
		5211: oled_colour = 16'b00000_000000_00000;
		5212: oled_colour = 16'b00000_000000_00000;
		5213: oled_colour = 16'b00000_000000_00000;
		5214: oled_colour = 16'b00000_000000_00000;
		5215: oled_colour = 16'b00000_000000_00000;
		5216: oled_colour = 16'b00000_000000_00000;
		5217: oled_colour = 16'b00000_000000_00000;
		5218: oled_colour = 16'b00000_000000_00000;
		5219: oled_colour = 16'b00000_000000_00000;
		5220: oled_colour = 16'b00000_000000_00000;
		5221: oled_colour = 16'b00000_000000_00000;
		5222: oled_colour = 16'b00000_000000_00000;
		5223: oled_colour = 16'b00000_000000_00000;
		5224: oled_colour = 16'b00000_000000_00000;
		5225: oled_colour = 16'b00000_000000_00000;
		5226: oled_colour = 16'b00000_000000_00000;
		5227: oled_colour = 16'b00000_000000_00000;
		5228: oled_colour = 16'b00000_000000_00000;
		5229: oled_colour = 16'b00000_000000_00000;
		5230: oled_colour = 16'b00000_000000_00000;
		5231: oled_colour = 16'b00000_000000_00000;
		5232: oled_colour = 16'b00000_000000_00000;
		5233: oled_colour = 16'b00000_000000_00000;
		5234: oled_colour = 16'b00000_000000_00000;
		5235: oled_colour = 16'b00000_000000_00000;
		5236: oled_colour = 16'b00000_000000_00000;
		5237: oled_colour = 16'b00000_000000_00000;
		5238: oled_colour = 16'b00000_000000_00000;
		5239: oled_colour = 16'b00000_000000_00000;
		5240: oled_colour = 16'b00000_000000_00000;
		5241: oled_colour = 16'b00000_000000_00000;
		5242: oled_colour = 16'b00000_000000_00000;
		5243: oled_colour = 16'b00000_000000_00000;
		5244: oled_colour = 16'b00000_000000_00000;
		5245: oled_colour = 16'b00000_000000_00000;
		5246: oled_colour = 16'b00000_000000_00000;
		5247: oled_colour = 16'b00000_000000_00000;
		5248: oled_colour = 16'b00000_000000_00000;
		5249: oled_colour = 16'b00000_000000_00000;
		5250: oled_colour = 16'b00000_000000_00000;
		5251: oled_colour = 16'b00000_000000_00000;
		5252: oled_colour = 16'b00000_000000_00000;
		5253: oled_colour = 16'b00000_000000_00000;
		5254: oled_colour = 16'b00000_000000_00000;
		5255: oled_colour = 16'b00000_000000_00000;
		5256: oled_colour = 16'b00000_000000_00000;
		5257: oled_colour = 16'b00000_000000_00000;
		5258: oled_colour = 16'b00000_000000_00000;
		5259: oled_colour = 16'b00000_000000_00000;
		5260: oled_colour = 16'b00000_000000_00000;
		5261: oled_colour = 16'b00000_000000_00000;
		5262: oled_colour = 16'b00000_000000_00000;
		5263: oled_colour = 16'b00000_000000_00000;
		5264: oled_colour = 16'b00000_000000_00000;
		5265: oled_colour = 16'b00000_000000_00000;
		5266: oled_colour = 16'b00000_000000_00000;
		5267: oled_colour = 16'b00000_000000_00000;
		5268: oled_colour = 16'b00000_000000_00000;
		5269: oled_colour = 16'b00000_000000_00000;
		5270: oled_colour = 16'b00000_000000_00000;
		5271: oled_colour = 16'b00000_000000_00000;
		5272: oled_colour = 16'b00000_000000_00000;
		5273: oled_colour = 16'b00000_000000_00000;
		5274: oled_colour = 16'b00000_000000_00000;
		5275: oled_colour = 16'b00000_000000_00000;
		5276: oled_colour = 16'b00000_000000_00000;
		5277: oled_colour = 16'b00000_000000_00000;
		5278: oled_colour = 16'b00000_000000_00000;
		5279: oled_colour = 16'b00000_000000_00000;
		5280: oled_colour = 16'b00000_000000_00000;
		5281: oled_colour = 16'b00000_000000_00000;
		5282: oled_colour = 16'b00000_000000_00000;
		5283: oled_colour = 16'b00000_000000_00000;
		5284: oled_colour = 16'b00000_000000_00000;
		5285: oled_colour = 16'b00000_000000_00000;
		5286: oled_colour = 16'b00000_000000_00000;
		5287: oled_colour = 16'b00000_000000_00000;
		5288: oled_colour = 16'b00000_000000_00000;
		5289: oled_colour = 16'b00000_000000_00000;
		5290: oled_colour = 16'b00000_000000_00000;
		5291: oled_colour = 16'b00000_000000_00000;
		5292: oled_colour = 16'b00000_000000_00000;
		5293: oled_colour = 16'b00000_000000_00000;
		5294: oled_colour = 16'b00000_000000_00000;
		5295: oled_colour = 16'b00000_000000_00000;
		5296: oled_colour = 16'b00000_000000_00000;
		5297: oled_colour = 16'b00000_000000_00000;
		5298: oled_colour = 16'b00000_000000_00000;
		5299: oled_colour = 16'b00000_000000_00000;
		5300: oled_colour = 16'b00000_000000_00000;
		5301: oled_colour = 16'b00000_000000_00000;
		5302: oled_colour = 16'b00000_000000_00000;
		5303: oled_colour = 16'b00000_000000_00000;
		5304: oled_colour = 16'b00000_000000_00000;
		5305: oled_colour = 16'b00000_000000_00000;
		5306: oled_colour = 16'b00000_000000_00000;
		5307: oled_colour = 16'b00000_000000_00000;
		5308: oled_colour = 16'b00000_000000_00000;
		5309: oled_colour = 16'b00000_000000_00000;
		5310: oled_colour = 16'b00000_000000_00000;
		5311: oled_colour = 16'b00000_000000_00000;
		5312: oled_colour = 16'b00000_000000_00000;
		5313: oled_colour = 16'b00000_000000_00000;
		5314: oled_colour = 16'b00000_000000_00000;
		5315: oled_colour = 16'b00000_000000_00000;
		5316: oled_colour = 16'b00000_000000_00000;
		5317: oled_colour = 16'b00000_000000_00000;
		5318: oled_colour = 16'b00000_000000_00000;
		5319: oled_colour = 16'b00000_000000_00000;
		5320: oled_colour = 16'b00000_000000_00000;
		5321: oled_colour = 16'b00000_000000_00000;
		5322: oled_colour = 16'b00000_000000_00000;
		5323: oled_colour = 16'b00000_000000_00000;
		5324: oled_colour = 16'b00000_000000_00000;
		5325: oled_colour = 16'b00000_000000_00000;
		5326: oled_colour = 16'b00000_000000_00000;
		5327: oled_colour = 16'b00000_000000_00000;
		5328: oled_colour = 16'b00000_000000_00000;
		5329: oled_colour = 16'b00000_000000_00000;
		5330: oled_colour = 16'b00000_000000_00000;
		5331: oled_colour = 16'b00000_000000_00000;
		5332: oled_colour = 16'b00000_000000_00000;
		5333: oled_colour = 16'b00000_000000_00000;
		5334: oled_colour = 16'b00000_000000_00000;
		5335: oled_colour = 16'b00000_000000_00000;
		5336: oled_colour = 16'b00000_000000_00000;
		5337: oled_colour = 16'b00000_000000_00000;
		5338: oled_colour = 16'b00000_000000_00000;
		5339: oled_colour = 16'b00000_000000_00000;
		5340: oled_colour = 16'b00000_000000_00000;
		5341: oled_colour = 16'b00000_000000_00000;
		5342: oled_colour = 16'b00000_000000_00000;
		5343: oled_colour = 16'b00000_000000_00000;
		5344: oled_colour = 16'b00000_000000_00000;
		5345: oled_colour = 16'b00000_000000_00000;
		5346: oled_colour = 16'b00000_000000_00000;
		5347: oled_colour = 16'b00000_000000_00000;
		5348: oled_colour = 16'b00000_000000_00000;
		5349: oled_colour = 16'b00000_000000_00000;
		5350: oled_colour = 16'b00000_000000_00000;
		5351: oled_colour = 16'b00000_000000_00000;
		5352: oled_colour = 16'b00000_000000_00000;
		5353: oled_colour = 16'b00000_000000_00000;
		5354: oled_colour = 16'b00000_000000_00000;
		5355: oled_colour = 16'b00000_000000_00000;
		5356: oled_colour = 16'b00000_000000_00000;
		5357: oled_colour = 16'b00000_000000_00000;
		5358: oled_colour = 16'b00000_000000_00000;
		5359: oled_colour = 16'b00000_000000_00000;
		5360: oled_colour = 16'b00000_000000_00000;
		5361: oled_colour = 16'b00000_000000_00000;
		5362: oled_colour = 16'b00000_000000_00000;
		5363: oled_colour = 16'b00000_000000_00000;
		5364: oled_colour = 16'b00000_000000_00000;
		5365: oled_colour = 16'b00000_000000_00000;
		5366: oled_colour = 16'b00000_000000_00000;
		5367: oled_colour = 16'b00000_000000_00000;
		5368: oled_colour = 16'b00000_000000_00000;
		5369: oled_colour = 16'b00000_000000_00000;
		5370: oled_colour = 16'b00000_000000_00000;
		5371: oled_colour = 16'b00000_000000_00000;
		5372: oled_colour = 16'b00000_000000_00000;
		5373: oled_colour = 16'b00000_000000_00000;
		5374: oled_colour = 16'b00000_000000_00000;
		5375: oled_colour = 16'b00000_000000_00000;
		5376: oled_colour = 16'b00000_000000_00000;
		5377: oled_colour = 16'b00000_000000_00000;
		5378: oled_colour = 16'b00000_000000_00000;
		5379: oled_colour = 16'b00000_000000_00000;
		5380: oled_colour = 16'b00000_000000_00000;
		5381: oled_colour = 16'b00000_000000_00000;
		5382: oled_colour = 16'b00000_000000_00000;
		5383: oled_colour = 16'b00000_000000_00000;
		5384: oled_colour = 16'b00000_000000_00000;
		5385: oled_colour = 16'b00000_000000_00000;
		5386: oled_colour = 16'b00000_000000_00000;
		5387: oled_colour = 16'b00000_000000_00000;
		5388: oled_colour = 16'b00000_000000_00000;
		5389: oled_colour = 16'b00000_000000_00000;
		5390: oled_colour = 16'b00000_000000_00000;
		5391: oled_colour = 16'b00000_000000_00000;
		5392: oled_colour = 16'b00000_000000_00000;
		5393: oled_colour = 16'b00000_000000_00000;
		5394: oled_colour = 16'b00000_000000_00000;
		5395: oled_colour = 16'b00000_000000_00000;
		5396: oled_colour = 16'b00000_000000_00000;
		5397: oled_colour = 16'b00000_000000_00000;
		5398: oled_colour = 16'b00000_000000_00000;
		5399: oled_colour = 16'b00000_000000_00000;
		5400: oled_colour = 16'b00000_000000_00000;
		5401: oled_colour = 16'b00000_000000_00000;
		5402: oled_colour = 16'b00000_000000_00000;
		5403: oled_colour = 16'b00000_000000_00000;
		5404: oled_colour = 16'b00000_000000_00000;
		5405: oled_colour = 16'b00000_000000_00000;
		5406: oled_colour = 16'b00000_000000_00000;
		5407: oled_colour = 16'b00000_000000_00000;
		5408: oled_colour = 16'b00000_000000_00000;
		5409: oled_colour = 16'b00000_000000_00000;
		5410: oled_colour = 16'b00000_000000_00000;
		5411: oled_colour = 16'b00000_000000_00000;
		5412: oled_colour = 16'b00000_000000_00000;
		5413: oled_colour = 16'b00000_000000_00000;
		5414: oled_colour = 16'b00000_000000_00000;
		5415: oled_colour = 16'b00000_000000_00000;
		5416: oled_colour = 16'b00000_000000_00000;
		5417: oled_colour = 16'b00000_000000_00000;
		5418: oled_colour = 16'b00000_000000_00000;
		5419: oled_colour = 16'b00000_000000_00000;
		5420: oled_colour = 16'b00000_000000_00000;
		5421: oled_colour = 16'b00000_000000_00000;
		5422: oled_colour = 16'b00000_000000_00000;
		5423: oled_colour = 16'b00000_000000_00000;
		5424: oled_colour = 16'b00000_000000_00000;
		5425: oled_colour = 16'b00000_000000_00000;
		5426: oled_colour = 16'b00000_000000_00000;
		5427: oled_colour = 16'b00000_000000_00000;
		5428: oled_colour = 16'b00000_000000_00000;
		5429: oled_colour = 16'b00000_000000_00000;
		5430: oled_colour = 16'b00000_000000_00000;
		5431: oled_colour = 16'b00000_000000_00000;
		5432: oled_colour = 16'b00000_000000_00000;
		5433: oled_colour = 16'b00000_000000_00000;
		5434: oled_colour = 16'b00000_000000_00000;
		5435: oled_colour = 16'b00000_000000_00000;
		5436: oled_colour = 16'b00000_000000_00000;
		5437: oled_colour = 16'b00000_000000_00000;
		5438: oled_colour = 16'b00000_000000_00000;
		5439: oled_colour = 16'b00000_000000_00000;
		5440: oled_colour = 16'b00000_000000_00000;
		5441: oled_colour = 16'b00000_000000_00000;
		5442: oled_colour = 16'b00000_000000_00000;
		5443: oled_colour = 16'b00000_000000_00000;
		5444: oled_colour = 16'b00000_000000_00000;
		5445: oled_colour = 16'b00000_000000_00000;
		5446: oled_colour = 16'b00000_000000_00000;
		5447: oled_colour = 16'b00000_000000_00000;
		5448: oled_colour = 16'b00000_000000_00000;
		5449: oled_colour = 16'b00000_000000_00000;
		5450: oled_colour = 16'b00000_000000_00000;
		5451: oled_colour = 16'b00000_000000_00000;
		5452: oled_colour = 16'b00000_000000_00000;
		5453: oled_colour = 16'b00000_000000_00000;
		5454: oled_colour = 16'b00000_000000_00000;
		5455: oled_colour = 16'b00000_000000_00000;
		5456: oled_colour = 16'b00000_000000_00000;
		5457: oled_colour = 16'b00000_000000_00000;
		5458: oled_colour = 16'b00000_000000_00000;
		5459: oled_colour = 16'b00000_000000_00000;
		5460: oled_colour = 16'b00000_000000_00000;
		5461: oled_colour = 16'b00000_000000_00000;
		5462: oled_colour = 16'b00000_000000_00000;
		5463: oled_colour = 16'b00000_000000_00000;
		5464: oled_colour = 16'b00000_000000_00000;
		5465: oled_colour = 16'b00000_000000_00000;
		5466: oled_colour = 16'b00000_000000_00000;
		5467: oled_colour = 16'b00000_000000_00000;
		5468: oled_colour = 16'b00000_000000_00000;
		5469: oled_colour = 16'b00000_000000_00000;
		5470: oled_colour = 16'b00000_000000_00000;
		5471: oled_colour = 16'b00000_000000_00000;
		5472: oled_colour = 16'b00000_000000_00000;
		5473: oled_colour = 16'b00000_000000_00000;
		5474: oled_colour = 16'b00000_000000_00000;
		5475: oled_colour = 16'b00000_000000_00000;
		5476: oled_colour = 16'b00000_000000_00000;
		5477: oled_colour = 16'b00000_000000_00000;
		5478: oled_colour = 16'b00000_000000_00000;
		5479: oled_colour = 16'b00000_000000_00000;
		5480: oled_colour = 16'b00000_000000_00000;
		5481: oled_colour = 16'b00000_000000_00000;
		5482: oled_colour = 16'b00000_000000_00000;
		5483: oled_colour = 16'b00000_000000_00000;
		5484: oled_colour = 16'b00000_000000_00000;
		5485: oled_colour = 16'b00000_000000_00000;
		5486: oled_colour = 16'b00000_000000_00000;
		5487: oled_colour = 16'b00000_000000_00000;
		5488: oled_colour = 16'b00000_000000_00000;
		5489: oled_colour = 16'b00000_000000_00000;
		5490: oled_colour = 16'b00000_000000_00000;
		5491: oled_colour = 16'b00000_000000_00000;
		5492: oled_colour = 16'b00000_000000_00000;
		5493: oled_colour = 16'b00000_000000_00000;
		5494: oled_colour = 16'b00000_000000_00000;
		5495: oled_colour = 16'b00000_000000_00000;
		5496: oled_colour = 16'b00000_000000_00000;
		5497: oled_colour = 16'b00000_000000_00000;
		5498: oled_colour = 16'b00000_000000_00000;
		5499: oled_colour = 16'b00000_000000_00000;
		5500: oled_colour = 16'b00000_000000_00000;
		5501: oled_colour = 16'b00000_000000_00000;
		5502: oled_colour = 16'b00000_000000_00000;
		5503: oled_colour = 16'b00000_000000_00000;
		5504: oled_colour = 16'b00000_000000_00000;
		5505: oled_colour = 16'b00000_000000_00000;
		5506: oled_colour = 16'b00000_000000_00000;
		5507: oled_colour = 16'b00000_000000_00000;
		5508: oled_colour = 16'b00000_000000_00000;
		5509: oled_colour = 16'b00000_000000_00000;
		5510: oled_colour = 16'b00000_000000_00000;
		5511: oled_colour = 16'b00000_000000_00000;
		5512: oled_colour = 16'b00000_000000_00000;
		5513: oled_colour = 16'b00000_000000_00000;
		5514: oled_colour = 16'b00000_000000_00000;
		5515: oled_colour = 16'b00000_000000_00000;
		5516: oled_colour = 16'b00000_000000_00000;
		5517: oled_colour = 16'b00000_000000_00000;
		5518: oled_colour = 16'b00000_000000_00000;
		5519: oled_colour = 16'b00000_000000_00000;
		5520: oled_colour = 16'b00000_000000_00000;
		5521: oled_colour = 16'b00000_000000_00000;
		5522: oled_colour = 16'b00000_000000_00000;
		5523: oled_colour = 16'b00000_000000_00000;
		5524: oled_colour = 16'b00000_000000_00000;
		5525: oled_colour = 16'b00000_000000_00000;
		5526: oled_colour = 16'b00000_000000_00000;
		5527: oled_colour = 16'b00000_000000_00000;
		5528: oled_colour = 16'b00000_000000_00000;
		5529: oled_colour = 16'b00000_000000_00000;
		5530: oled_colour = 16'b00000_000000_00000;
		5531: oled_colour = 16'b00000_000000_00000;
		5532: oled_colour = 16'b00000_000000_00000;
		5533: oled_colour = 16'b00000_000000_00000;
		5534: oled_colour = 16'b00000_000000_00000;
		5535: oled_colour = 16'b00000_000000_00000;
		5536: oled_colour = 16'b00000_000000_00000;
		5537: oled_colour = 16'b00000_000000_00000;
		5538: oled_colour = 16'b00000_000000_00000;
		5539: oled_colour = 16'b00000_000000_00000;
		5540: oled_colour = 16'b00000_000000_00000;
		5541: oled_colour = 16'b00000_000000_00000;
		5542: oled_colour = 16'b00000_000000_00000;
		5543: oled_colour = 16'b00000_000000_00000;
		5544: oled_colour = 16'b00000_000000_00000;
		5545: oled_colour = 16'b00000_000000_00000;
		5546: oled_colour = 16'b00000_000000_00000;
		5547: oled_colour = 16'b00000_000000_00000;
		5548: oled_colour = 16'b00000_000000_00000;
		5549: oled_colour = 16'b00000_000000_00000;
		5550: oled_colour = 16'b00000_000000_00000;
		5551: oled_colour = 16'b00000_000000_00000;
		5552: oled_colour = 16'b00000_000000_00000;
		5553: oled_colour = 16'b00000_000000_00000;
		5554: oled_colour = 16'b00000_000000_00000;
		5555: oled_colour = 16'b00000_000000_00000;
		5556: oled_colour = 16'b00000_000000_00000;
		5557: oled_colour = 16'b00000_000000_00000;
		5558: oled_colour = 16'b00000_000000_00000;
		5559: oled_colour = 16'b00000_000000_00000;
		5560: oled_colour = 16'b00000_000000_00000;
		5561: oled_colour = 16'b00000_000000_00000;
		5562: oled_colour = 16'b00000_000000_00000;
		5563: oled_colour = 16'b00000_000000_00000;
		5564: oled_colour = 16'b00000_000000_00000;
		5565: oled_colour = 16'b00000_000000_00000;
		5566: oled_colour = 16'b00000_000000_00000;
		5567: oled_colour = 16'b00000_000000_00000;
		5568: oled_colour = 16'b00000_000000_00000;
		5569: oled_colour = 16'b00000_000000_00000;
		5570: oled_colour = 16'b00000_000000_00000;
		5571: oled_colour = 16'b00000_000000_00000;
		5572: oled_colour = 16'b00000_000000_00000;
		5573: oled_colour = 16'b00000_000000_00000;
		5574: oled_colour = 16'b00000_000000_00000;
		5575: oled_colour = 16'b00000_000000_00000;
		5576: oled_colour = 16'b00000_000000_00000;
		5577: oled_colour = 16'b00000_000000_00000;
		5578: oled_colour = 16'b00000_000000_00000;
		5579: oled_colour = 16'b00000_000000_00000;
		5580: oled_colour = 16'b00000_000000_00000;
		5581: oled_colour = 16'b00000_000000_00000;
		5582: oled_colour = 16'b00000_000000_00000;
		5583: oled_colour = 16'b00000_000000_00000;
		5584: oled_colour = 16'b00000_000000_00000;
		5585: oled_colour = 16'b00000_000000_00000;
		5586: oled_colour = 16'b00000_000000_00000;
		5587: oled_colour = 16'b00000_000000_00000;
		5588: oled_colour = 16'b00000_000000_00000;
		5589: oled_colour = 16'b00000_000000_00000;
		5590: oled_colour = 16'b00000_000000_00000;
		5591: oled_colour = 16'b00000_000000_00000;
		5592: oled_colour = 16'b00000_000000_00000;
		5593: oled_colour = 16'b00000_000000_00000;
		5594: oled_colour = 16'b00000_000000_00000;
		5595: oled_colour = 16'b00000_000000_00000;
		5596: oled_colour = 16'b00000_000000_00000;
		5597: oled_colour = 16'b00000_000000_00000;
		5598: oled_colour = 16'b00000_000000_00000;
		5599: oled_colour = 16'b00000_000000_00000;
		5600: oled_colour = 16'b00000_000000_00000;
		5601: oled_colour = 16'b00000_000000_00000;
		5602: oled_colour = 16'b00000_000000_00000;
		5603: oled_colour = 16'b00000_000000_00000;
		5604: oled_colour = 16'b00000_000000_00000;
		5605: oled_colour = 16'b00000_000000_00000;
		5606: oled_colour = 16'b00000_000000_00000;
		5607: oled_colour = 16'b00000_000000_00000;
		5608: oled_colour = 16'b00000_000000_00000;
		5609: oled_colour = 16'b00000_000000_00000;
		5610: oled_colour = 16'b00000_000000_00000;
		5611: oled_colour = 16'b00000_000000_00000;
		5612: oled_colour = 16'b00000_000000_00000;
		5613: oled_colour = 16'b00000_000000_00000;
		5614: oled_colour = 16'b00000_000000_00000;
		5615: oled_colour = 16'b00000_000000_00000;
		5616: oled_colour = 16'b00000_000000_00000;
		5617: oled_colour = 16'b00000_000000_00000;
		5618: oled_colour = 16'b00000_000000_00000;
		5619: oled_colour = 16'b00000_000000_00000;
		5620: oled_colour = 16'b00000_000000_00000;
		5621: oled_colour = 16'b00000_000000_00000;
		5622: oled_colour = 16'b00000_000000_00000;
		5623: oled_colour = 16'b00000_000000_00000;
		5624: oled_colour = 16'b00000_000000_00000;
		5625: oled_colour = 16'b00000_000000_00000;
		5626: oled_colour = 16'b00000_000000_00000;
		5627: oled_colour = 16'b00000_000000_00000;
		5628: oled_colour = 16'b00000_000000_00000;
		5629: oled_colour = 16'b00000_000000_00000;
		5630: oled_colour = 16'b00000_000000_00000;
		5631: oled_colour = 16'b00000_000000_00000;
		5632: oled_colour = 16'b00000_000000_00000;
		5633: oled_colour = 16'b00000_000000_00000;
		5634: oled_colour = 16'b00000_000000_00000;
		5635: oled_colour = 16'b00000_000000_00000;
		5636: oled_colour = 16'b00000_000000_00000;
		5637: oled_colour = 16'b00000_000000_00000;
		5638: oled_colour = 16'b00000_000000_00000;
		5639: oled_colour = 16'b00000_000000_00000;
		5640: oled_colour = 16'b00000_000000_00000;
		5641: oled_colour = 16'b00000_000000_00000;
		5642: oled_colour = 16'b00000_000000_00000;
		5643: oled_colour = 16'b00000_000000_00000;
		5644: oled_colour = 16'b00000_000000_00000;
		5645: oled_colour = 16'b00000_000000_00000;
		5646: oled_colour = 16'b00000_000000_00000;
		5647: oled_colour = 16'b00000_000000_00000;
		5648: oled_colour = 16'b00000_000000_00000;
		5649: oled_colour = 16'b00000_000000_00000;
		5650: oled_colour = 16'b00000_000000_00000;
		5651: oled_colour = 16'b00000_000000_00000;
		5652: oled_colour = 16'b00000_000000_00000;
		5653: oled_colour = 16'b00000_000000_00000;
		5654: oled_colour = 16'b00000_000000_00000;
		5655: oled_colour = 16'b00000_000000_00000;
		5656: oled_colour = 16'b00000_000000_00000;
		5657: oled_colour = 16'b00000_000000_00000;
		5658: oled_colour = 16'b00000_000000_00000;
		5659: oled_colour = 16'b00000_000000_00000;
		5660: oled_colour = 16'b00000_000000_00000;
		5661: oled_colour = 16'b00000_000000_00000;
		5662: oled_colour = 16'b00000_000000_00000;
		5663: oled_colour = 16'b00000_000000_00000;
		5664: oled_colour = 16'b00000_000000_00000;
		5665: oled_colour = 16'b00000_000000_00000;
		5666: oled_colour = 16'b00000_000000_00000;
		5667: oled_colour = 16'b00000_000000_00000;
		5668: oled_colour = 16'b00000_000000_00000;
		5669: oled_colour = 16'b00000_000000_00000;
		5670: oled_colour = 16'b00000_000000_00000;
		5671: oled_colour = 16'b00000_000000_00000;
		5672: oled_colour = 16'b00000_000000_00000;
		5673: oled_colour = 16'b00000_000000_00000;
		5674: oled_colour = 16'b00000_000000_00000;
		5675: oled_colour = 16'b00000_000000_00000;
		5676: oled_colour = 16'b00000_000000_00000;
		5677: oled_colour = 16'b00000_000000_00000;
		5678: oled_colour = 16'b00000_000000_00000;
		5679: oled_colour = 16'b00000_000000_00000;
		5680: oled_colour = 16'b00000_000000_00000;
		5681: oled_colour = 16'b00000_000000_00000;
		5682: oled_colour = 16'b00000_000000_00000;
		5683: oled_colour = 16'b00000_000000_00000;
		5684: oled_colour = 16'b00000_000000_00000;
		5685: oled_colour = 16'b00000_000000_00000;
		5686: oled_colour = 16'b00000_000000_00000;
		5687: oled_colour = 16'b00000_000000_00000;
		5688: oled_colour = 16'b00000_000000_00000;
		5689: oled_colour = 16'b00000_000000_00000;
		5690: oled_colour = 16'b00000_000000_00000;
		5691: oled_colour = 16'b00000_000000_00000;
		5692: oled_colour = 16'b00000_000000_00000;
		5693: oled_colour = 16'b00000_000000_00000;
		5694: oled_colour = 16'b00000_000000_00000;
		5695: oled_colour = 16'b00000_000000_00000;
		5696: oled_colour = 16'b00000_000000_00000;
		5697: oled_colour = 16'b00000_000000_00000;
		5698: oled_colour = 16'b00000_000000_00000;
		5699: oled_colour = 16'b00000_000000_00000;
		5700: oled_colour = 16'b00000_000000_00000;
		5701: oled_colour = 16'b00000_000000_00000;
		5702: oled_colour = 16'b00000_000000_00000;
		5703: oled_colour = 16'b00000_000000_00000;
		5704: oled_colour = 16'b00000_000000_00000;
		5705: oled_colour = 16'b00000_000000_00000;
		5706: oled_colour = 16'b00000_000000_00000;
		5707: oled_colour = 16'b00000_000000_00000;
		5708: oled_colour = 16'b00000_000000_00000;
		5709: oled_colour = 16'b00000_000000_00000;
		5710: oled_colour = 16'b00000_000000_00000;
		5711: oled_colour = 16'b00000_000000_00000;
		5712: oled_colour = 16'b00000_000000_00000;
		5713: oled_colour = 16'b00000_000000_00000;
		5714: oled_colour = 16'b00000_000000_00000;
		5715: oled_colour = 16'b00000_000000_00000;
		5716: oled_colour = 16'b00000_000000_00000;
		5717: oled_colour = 16'b00000_000000_00000;
		5718: oled_colour = 16'b00000_000000_00000;
		5719: oled_colour = 16'b00000_000000_00000;
		5720: oled_colour = 16'b00000_000000_00000;
		5721: oled_colour = 16'b00000_000000_00000;
		5722: oled_colour = 16'b00000_000000_00000;
		5723: oled_colour = 16'b00000_000000_00000;
		5724: oled_colour = 16'b00000_000000_00000;
		5725: oled_colour = 16'b00000_000000_00000;
		5726: oled_colour = 16'b00000_000000_00000;
		5727: oled_colour = 16'b00000_000000_00000;
		5728: oled_colour = 16'b00000_000000_00000;
		5729: oled_colour = 16'b00000_000000_00000;
		5730: oled_colour = 16'b00000_000000_00000;
		5731: oled_colour = 16'b00000_000000_00000;
		5732: oled_colour = 16'b00000_000000_00000;
		5733: oled_colour = 16'b00000_000000_00000;
		5734: oled_colour = 16'b00000_000000_00000;
		5735: oled_colour = 16'b00000_000000_00000;
		5736: oled_colour = 16'b00000_000000_00000;
		5737: oled_colour = 16'b00000_000000_00000;
		5738: oled_colour = 16'b00000_000000_00000;
		5739: oled_colour = 16'b00000_000000_00000;
		5740: oled_colour = 16'b00000_000000_00000;
		5741: oled_colour = 16'b00000_000000_00000;
		5742: oled_colour = 16'b00000_000000_00000;
		5743: oled_colour = 16'b00000_000000_00000;
		5744: oled_colour = 16'b00000_000000_00000;
		5745: oled_colour = 16'b00000_000000_00000;
		5746: oled_colour = 16'b00000_000000_00000;
		5747: oled_colour = 16'b00000_000000_00000;
		5748: oled_colour = 16'b00000_000000_00000;
		5749: oled_colour = 16'b00000_000000_00000;
		5750: oled_colour = 16'b00000_000000_00000;
		5751: oled_colour = 16'b00000_000000_00000;
		5752: oled_colour = 16'b00000_000000_00000;
		5753: oled_colour = 16'b00000_000000_00000;
		5754: oled_colour = 16'b00000_000000_00000;
		5755: oled_colour = 16'b00000_000000_00000;
		5756: oled_colour = 16'b00000_000000_00000;
		5757: oled_colour = 16'b00000_000000_00000;
		5758: oled_colour = 16'b00000_000000_00000;
		5759: oled_colour = 16'b00000_000000_00000;
		5760: oled_colour = 16'b00000_000000_00000;
		5761: oled_colour = 16'b00000_000000_00000;
		5762: oled_colour = 16'b00000_000000_00000;
		5763: oled_colour = 16'b00000_000000_00000;
		5764: oled_colour = 16'b00000_000000_00000;
		5765: oled_colour = 16'b00000_000000_00000;
		5766: oled_colour = 16'b00000_000000_00000;
		5767: oled_colour = 16'b00000_000000_00000;
		5768: oled_colour = 16'b00000_000000_00000;
		5769: oled_colour = 16'b00000_000000_00000;
		5770: oled_colour = 16'b00000_000000_00000;
		5771: oled_colour = 16'b00000_000000_00000;
		5772: oled_colour = 16'b00000_000000_00000;
		5773: oled_colour = 16'b00000_000000_00000;
		5774: oled_colour = 16'b00000_000000_00000;
		5775: oled_colour = 16'b00000_000000_00000;
		5776: oled_colour = 16'b00000_000000_00000;
		5777: oled_colour = 16'b00000_000000_00000;
		5778: oled_colour = 16'b00000_000000_00000;
		5779: oled_colour = 16'b00000_000000_00000;
		5780: oled_colour = 16'b00000_000000_00000;
		5781: oled_colour = 16'b00000_000000_00000;
		5782: oled_colour = 16'b00000_000000_00000;
		5783: oled_colour = 16'b00000_000000_00000;
		5784: oled_colour = 16'b00000_000000_00000;
		5785: oled_colour = 16'b00000_000000_00000;
		5786: oled_colour = 16'b00000_000000_00000;
		5787: oled_colour = 16'b00000_000000_00000;
		5788: oled_colour = 16'b00000_000000_00000;
		5789: oled_colour = 16'b00000_000000_00000;
		5790: oled_colour = 16'b00000_000000_00000;
		5791: oled_colour = 16'b00000_000000_00000;
		5792: oled_colour = 16'b00000_000000_00000;
		5793: oled_colour = 16'b00000_000000_00000;
		5794: oled_colour = 16'b00000_000000_00000;
		5795: oled_colour = 16'b00000_000000_00000;
		5796: oled_colour = 16'b00000_000000_00000;
		5797: oled_colour = 16'b00000_000000_00000;
		5798: oled_colour = 16'b00000_000000_00000;
		5799: oled_colour = 16'b00000_000000_00000;
		5800: oled_colour = 16'b00000_000000_00000;
		5801: oled_colour = 16'b00000_000000_00000;
		5802: oled_colour = 16'b00000_000000_00000;
		5803: oled_colour = 16'b00000_000000_00000;
		5804: oled_colour = 16'b00000_000000_00000;
		5805: oled_colour = 16'b00000_000000_00000;
		5806: oled_colour = 16'b00000_000000_00000;
		5807: oled_colour = 16'b00000_000000_00000;
		5808: oled_colour = 16'b00000_000000_00000;
		5809: oled_colour = 16'b00000_000000_00000;
		5810: oled_colour = 16'b00000_000000_00000;
		5811: oled_colour = 16'b00000_000000_00000;
		5812: oled_colour = 16'b00000_000000_00000;
		5813: oled_colour = 16'b00000_000000_00000;
		5814: oled_colour = 16'b00000_000000_00000;
		5815: oled_colour = 16'b00000_000000_00000;
		5816: oled_colour = 16'b00000_000000_00000;
		5817: oled_colour = 16'b00000_000000_00000;
		5818: oled_colour = 16'b00000_000000_00000;
		5819: oled_colour = 16'b00000_000000_00000;
		5820: oled_colour = 16'b00000_000000_00000;
		5821: oled_colour = 16'b00000_000000_00000;
		5822: oled_colour = 16'b00000_000000_00000;
		5823: oled_colour = 16'b00000_000000_00000;
		5824: oled_colour = 16'b00000_000000_00000;
		5825: oled_colour = 16'b00000_000000_00000;
		5826: oled_colour = 16'b00000_000000_00000;
		5827: oled_colour = 16'b00000_000000_00000;
		5828: oled_colour = 16'b00000_000000_00000;
		5829: oled_colour = 16'b00000_000000_00000;
		5830: oled_colour = 16'b00000_000000_00000;
		5831: oled_colour = 16'b00000_000000_00000;
		5832: oled_colour = 16'b00000_000000_00000;
		5833: oled_colour = 16'b00000_000000_00000;
		5834: oled_colour = 16'b00000_000000_00000;
		5835: oled_colour = 16'b00000_000000_00000;
		5836: oled_colour = 16'b00000_000000_00000;
		5837: oled_colour = 16'b00000_000000_00000;
		5838: oled_colour = 16'b00000_000000_00000;
		5839: oled_colour = 16'b00000_000000_00000;
		5840: oled_colour = 16'b00000_000000_00000;
		5841: oled_colour = 16'b00000_000000_00000;
		5842: oled_colour = 16'b00000_000000_00000;
		5843: oled_colour = 16'b00000_000000_00000;
		5844: oled_colour = 16'b00000_000000_00000;
		5845: oled_colour = 16'b00000_000000_00000;
		5846: oled_colour = 16'b00000_000000_00000;
		5847: oled_colour = 16'b00000_000000_00000;
		5848: oled_colour = 16'b00000_000000_00000;
		5849: oled_colour = 16'b00000_000000_00000;
		5850: oled_colour = 16'b00000_000000_00000;
		5851: oled_colour = 16'b00000_000000_00000;
		5852: oled_colour = 16'b00000_000000_00000;
		5853: oled_colour = 16'b00000_000000_00000;
		5854: oled_colour = 16'b00000_000000_00000;
		5855: oled_colour = 16'b00000_000000_00000;
		5856: oled_colour = 16'b00000_000000_00000;
		5857: oled_colour = 16'b00000_000000_00000;
		5858: oled_colour = 16'b00000_000000_00000;
		5859: oled_colour = 16'b00000_000000_00000;
		5860: oled_colour = 16'b00000_000000_00000;
		5861: oled_colour = 16'b00000_000000_00000;
		5862: oled_colour = 16'b00000_000000_00000;
		5863: oled_colour = 16'b00000_000000_00000;
		5864: oled_colour = 16'b00000_000000_00000;
		5865: oled_colour = 16'b00000_000000_00000;
		5866: oled_colour = 16'b00000_000000_00000;
		5867: oled_colour = 16'b00000_000000_00000;
		5868: oled_colour = 16'b00000_000000_00000;
		5869: oled_colour = 16'b00000_000000_00000;
		5870: oled_colour = 16'b00000_000000_00000;
		5871: oled_colour = 16'b00000_000000_00000;
		5872: oled_colour = 16'b00000_000000_00000;
		5873: oled_colour = 16'b00000_000000_00000;
		5874: oled_colour = 16'b00000_000000_00000;
		5875: oled_colour = 16'b00000_000000_00000;
		5876: oled_colour = 16'b00000_000000_00000;
		5877: oled_colour = 16'b00000_000000_00000;
		5878: oled_colour = 16'b00000_000000_00000;
		5879: oled_colour = 16'b00000_000000_00000;
		5880: oled_colour = 16'b00000_000000_00000;
		5881: oled_colour = 16'b00000_000000_00000;
		5882: oled_colour = 16'b00000_000000_00000;
		5883: oled_colour = 16'b00000_000000_00000;
		5884: oled_colour = 16'b00000_000000_00000;
		5885: oled_colour = 16'b00000_000000_00000;
		5886: oled_colour = 16'b00000_000000_00000;
		5887: oled_colour = 16'b00000_000000_00000;
		5888: oled_colour = 16'b00000_000000_00000;
		5889: oled_colour = 16'b00000_000000_00000;
		5890: oled_colour = 16'b00000_000000_00000;
		5891: oled_colour = 16'b00000_000000_00000;
		5892: oled_colour = 16'b00000_000000_00000;
		5893: oled_colour = 16'b00000_000000_00000;
		5894: oled_colour = 16'b00000_000000_00000;
		5895: oled_colour = 16'b00000_000000_00000;
		5896: oled_colour = 16'b00000_000000_00000;
		5897: oled_colour = 16'b00000_000000_00000;
		5898: oled_colour = 16'b00000_000000_00000;
		5899: oled_colour = 16'b00000_000000_00000;
		5900: oled_colour = 16'b00000_000000_00000;
		5901: oled_colour = 16'b00000_000000_00000;
		5902: oled_colour = 16'b00000_000000_00000;
		5903: oled_colour = 16'b00000_000000_00000;
		5904: oled_colour = 16'b00000_000000_00000;
		5905: oled_colour = 16'b00000_000000_00000;
		5906: oled_colour = 16'b00000_000000_00000;
		5907: oled_colour = 16'b00000_000000_00000;
		5908: oled_colour = 16'b00000_000000_00000;
		5909: oled_colour = 16'b00000_000000_00000;
		5910: oled_colour = 16'b00000_000000_00000;
		5911: oled_colour = 16'b00000_000000_00000;
		5912: oled_colour = 16'b00000_000000_00000;
		5913: oled_colour = 16'b00000_000000_00000;
		5914: oled_colour = 16'b00000_000000_00000;
		5915: oled_colour = 16'b00000_000000_00000;
		5916: oled_colour = 16'b00000_000000_00000;
		5917: oled_colour = 16'b00000_000000_00000;
		5918: oled_colour = 16'b00000_000000_00000;
		5919: oled_colour = 16'b00000_000000_00000;
		5920: oled_colour = 16'b00000_000000_00000;
		5921: oled_colour = 16'b00000_000000_00000;
		5922: oled_colour = 16'b00000_000000_00000;
		5923: oled_colour = 16'b00000_000000_00000;
		5924: oled_colour = 16'b00000_000000_00000;
		5925: oled_colour = 16'b00000_000000_00000;
		5926: oled_colour = 16'b00000_000000_00000;
		5927: oled_colour = 16'b00000_000000_00000;
		5928: oled_colour = 16'b00000_000000_00000;
		5929: oled_colour = 16'b00000_000000_00000;
		5930: oled_colour = 16'b00000_000000_00000;
		5931: oled_colour = 16'b00000_000000_00000;
		5932: oled_colour = 16'b00000_000000_00000;
		5933: oled_colour = 16'b00000_000000_00000;
		5934: oled_colour = 16'b00000_000000_00000;
		5935: oled_colour = 16'b00000_000000_00000;
		5936: oled_colour = 16'b00000_000000_00000;
		5937: oled_colour = 16'b00000_000000_00000;
		5938: oled_colour = 16'b00000_000000_00000;
		5939: oled_colour = 16'b00000_000000_00000;
		5940: oled_colour = 16'b00000_000000_00000;
		5941: oled_colour = 16'b00000_000000_00000;
		5942: oled_colour = 16'b00000_000000_00000;
		5943: oled_colour = 16'b00000_000000_00000;
		5944: oled_colour = 16'b00000_000000_00000;
		5945: oled_colour = 16'b00000_000000_00000;
		5946: oled_colour = 16'b00000_000000_00000;
		5947: oled_colour = 16'b00000_000000_00000;
		5948: oled_colour = 16'b00000_000000_00000;
		5949: oled_colour = 16'b00000_000000_00000;
		5950: oled_colour = 16'b00000_000000_00000;
		5951: oled_colour = 16'b00000_000000_00000;
		5952: oled_colour = 16'b00000_000000_00000;
		5953: oled_colour = 16'b00000_000000_00000;
		5954: oled_colour = 16'b00000_000000_00000;
		5955: oled_colour = 16'b00000_000000_00000;
		5956: oled_colour = 16'b00000_000000_00000;
		5957: oled_colour = 16'b00000_000000_00000;
		5958: oled_colour = 16'b00000_000000_00000;
		5959: oled_colour = 16'b00000_000000_00000;
		5960: oled_colour = 16'b00000_000000_00000;
		5961: oled_colour = 16'b00000_000000_00000;
		5962: oled_colour = 16'b00000_000000_00000;
		5963: oled_colour = 16'b00000_000000_00000;
		5964: oled_colour = 16'b00000_000000_00000;
		5965: oled_colour = 16'b00000_000000_00000;
		5966: oled_colour = 16'b00000_000000_00000;
		5967: oled_colour = 16'b00000_000000_00000;
		5968: oled_colour = 16'b00000_000000_00000;
		5969: oled_colour = 16'b00000_000000_00000;
		5970: oled_colour = 16'b00000_000000_00000;
		5971: oled_colour = 16'b00000_000000_00000;
		5972: oled_colour = 16'b00000_000000_00000;
		5973: oled_colour = 16'b00000_000000_00000;
		5974: oled_colour = 16'b00000_000000_00000;
		5975: oled_colour = 16'b00000_000000_00000;
		5976: oled_colour = 16'b00000_000000_00000;
		5977: oled_colour = 16'b00000_000000_00000;
		5978: oled_colour = 16'b00000_000000_00000;
		5979: oled_colour = 16'b00000_000000_00000;
		5980: oled_colour = 16'b00000_000000_00000;
		5981: oled_colour = 16'b00000_000000_00000;
		5982: oled_colour = 16'b00000_000000_00000;
		5983: oled_colour = 16'b00000_000000_00000;
		5984: oled_colour = 16'b00000_000000_00000;
		5985: oled_colour = 16'b00000_000000_00000;
		5986: oled_colour = 16'b00000_000000_00000;
		5987: oled_colour = 16'b00000_000000_00000;
		5988: oled_colour = 16'b00000_000000_00000;
		5989: oled_colour = 16'b00000_000000_00000;
		5990: oled_colour = 16'b00000_000000_00000;
		5991: oled_colour = 16'b00000_000000_00000;
		5992: oled_colour = 16'b00000_000000_00000;
		5993: oled_colour = 16'b00000_000000_00000;
		5994: oled_colour = 16'b00000_000000_00000;
		5995: oled_colour = 16'b00000_000000_00000;
		5996: oled_colour = 16'b00000_000000_00000;
		5997: oled_colour = 16'b00000_000000_00000;
		5998: oled_colour = 16'b00000_000000_00000;
		5999: oled_colour = 16'b00000_000000_00000;
		6000: oled_colour = 16'b00000_000000_00000;
		6001: oled_colour = 16'b00000_000000_00000;
		6002: oled_colour = 16'b00000_000000_00000;
		6003: oled_colour = 16'b00000_000000_00000;
		6004: oled_colour = 16'b00000_000000_00000;
		6005: oled_colour = 16'b00000_000000_00000;
		6006: oled_colour = 16'b00000_000000_00000;
		6007: oled_colour = 16'b00000_000000_00000;
		6008: oled_colour = 16'b00000_000000_00000;
		6009: oled_colour = 16'b00000_000000_00000;
		6010: oled_colour = 16'b00000_000000_00000;
		6011: oled_colour = 16'b00000_000000_00000;
		6012: oled_colour = 16'b00000_000000_00000;
		6013: oled_colour = 16'b00000_000000_00000;
		6014: oled_colour = 16'b00000_000000_00000;
		6015: oled_colour = 16'b00000_000000_00000;
		6016: oled_colour = 16'b00000_000000_00000;
		6017: oled_colour = 16'b00000_000000_00000;
		6018: oled_colour = 16'b00000_000000_00000;
		6019: oled_colour = 16'b00000_000000_00000;
		6020: oled_colour = 16'b00000_000000_00000;
		6021: oled_colour = 16'b00000_000000_00000;
		6022: oled_colour = 16'b00000_000000_00000;
		6023: oled_colour = 16'b00000_000000_00000;
		6024: oled_colour = 16'b00000_000000_00000;
		6025: oled_colour = 16'b00000_000000_00000;
		6026: oled_colour = 16'b00000_000000_00000;
		6027: oled_colour = 16'b00000_000000_00000;
		6028: oled_colour = 16'b00000_000000_00000;
		6029: oled_colour = 16'b00000_000000_00000;
		6030: oled_colour = 16'b00000_000000_00000;
		6031: oled_colour = 16'b00000_000000_00000;
		6032: oled_colour = 16'b00000_000000_00000;
		6033: oled_colour = 16'b00000_000000_00000;
		6034: oled_colour = 16'b00000_000000_00000;
		6035: oled_colour = 16'b00000_000000_00000;
		6036: oled_colour = 16'b00000_000000_00000;
		6037: oled_colour = 16'b00000_000000_00000;
		6038: oled_colour = 16'b00000_000000_00000;
		6039: oled_colour = 16'b00000_000000_00000;
		6040: oled_colour = 16'b00000_000000_00000;
		6041: oled_colour = 16'b00000_000000_00000;
		6042: oled_colour = 16'b00000_000000_00000;
		6043: oled_colour = 16'b00000_000000_00000;
		6044: oled_colour = 16'b00000_000000_00000;
		6045: oled_colour = 16'b00000_000000_00000;
		6046: oled_colour = 16'b00000_000000_00000;
		6047: oled_colour = 16'b00000_000000_00000;
		6048: oled_colour = 16'b00000_000000_00000;
		6049: oled_colour = 16'b00000_000000_00000;
		6050: oled_colour = 16'b00000_000000_00000;
		6051: oled_colour = 16'b00000_000000_00000;
		6052: oled_colour = 16'b00000_000000_00000;
		6053: oled_colour = 16'b00000_000000_00000;
		6054: oled_colour = 16'b00000_000000_00000;
		6055: oled_colour = 16'b00000_000000_00000;
		6056: oled_colour = 16'b00000_000000_00000;
		6057: oled_colour = 16'b00000_000000_00000;
		6058: oled_colour = 16'b00000_000000_00000;
		6059: oled_colour = 16'b00000_000000_00000;
		6060: oled_colour = 16'b00000_000000_00000;
		6061: oled_colour = 16'b00000_000000_00000;
		6062: oled_colour = 16'b00000_000000_00000;
		6063: oled_colour = 16'b00000_000000_00000;
		6064: oled_colour = 16'b00000_000000_00000;
		6065: oled_colour = 16'b00000_000000_00000;
		6066: oled_colour = 16'b00000_000000_00000;
		6067: oled_colour = 16'b00000_000000_00000;
		6068: oled_colour = 16'b00000_000000_00000;
		6069: oled_colour = 16'b00000_000000_00000;
		6070: oled_colour = 16'b00000_000000_00000;
		6071: oled_colour = 16'b00000_000000_00000;
		6072: oled_colour = 16'b00000_000000_00000;
		6073: oled_colour = 16'b00000_000000_00000;
		6074: oled_colour = 16'b00000_000000_00000;
		6075: oled_colour = 16'b00000_000000_00000;
		6076: oled_colour = 16'b00000_000000_00000;
		6077: oled_colour = 16'b00000_000000_00000;
		6078: oled_colour = 16'b00000_000000_00000;
		6079: oled_colour = 16'b00000_000000_00000;
		6080: oled_colour = 16'b00000_000000_00000;
		6081: oled_colour = 16'b00000_000000_00000;
		6082: oled_colour = 16'b00000_000000_00000;
		6083: oled_colour = 16'b00000_000000_00000;
		6084: oled_colour = 16'b00000_000000_00000;
		6085: oled_colour = 16'b00000_000000_00000;
		6086: oled_colour = 16'b00000_000000_00000;
		6087: oled_colour = 16'b00000_000000_00000;
		6088: oled_colour = 16'b00000_000000_00000;
		6089: oled_colour = 16'b00000_000000_00000;
		6090: oled_colour = 16'b00000_000000_00000;
		6091: oled_colour = 16'b00000_000000_00000;
		6092: oled_colour = 16'b00000_000000_00000;
		6093: oled_colour = 16'b00000_000000_00000;
		6094: oled_colour = 16'b00000_000000_00000;
		6095: oled_colour = 16'b00000_000000_00000;
		6096: oled_colour = 16'b00000_000000_00000;
		6097: oled_colour = 16'b00000_000000_00000;
		6098: oled_colour = 16'b00000_000000_00000;
		6099: oled_colour = 16'b00000_000000_00000;
		6100: oled_colour = 16'b00000_000000_00000;
		6101: oled_colour = 16'b00000_000000_00000;
		6102: oled_colour = 16'b00000_000000_00000;
		6103: oled_colour = 16'b00000_000000_00000;
		6104: oled_colour = 16'b00000_000000_00000;
		6105: oled_colour = 16'b00000_000000_00000;
		6106: oled_colour = 16'b00000_000000_00000;
		6107: oled_colour = 16'b00000_000000_00000;
		6108: oled_colour = 16'b00000_000000_00000;
		6109: oled_colour = 16'b00000_000000_00000;
		6110: oled_colour = 16'b00000_000000_00000;
		6111: oled_colour = 16'b00000_000000_00000;
		6112: oled_colour = 16'b00000_000000_00000;
		6113: oled_colour = 16'b00000_000000_00000;
		6114: oled_colour = 16'b00000_000000_00000;
		6115: oled_colour = 16'b00000_000000_00000;
		6116: oled_colour = 16'b00000_000000_00000;
		6117: oled_colour = 16'b00000_000000_00000;
		6118: oled_colour = 16'b00000_000000_00000;
		6119: oled_colour = 16'b00000_000000_00000;
		6120: oled_colour = 16'b00000_000000_00000;
		6121: oled_colour = 16'b00000_000000_00000;
		6122: oled_colour = 16'b00000_000000_00000;
		6123: oled_colour = 16'b00000_000000_00000;
		6124: oled_colour = 16'b00000_000000_00000;
		6125: oled_colour = 16'b00000_000000_00000;
		6126: oled_colour = 16'b00000_000000_00000;
		6127: oled_colour = 16'b00000_000000_00000;
		6128: oled_colour = 16'b00000_000000_00000;
		6129: oled_colour = 16'b00000_000000_00000;
		6130: oled_colour = 16'b00000_000000_00000;
		6131: oled_colour = 16'b00000_000000_00000;
		6132: oled_colour = 16'b00000_000000_00000;
		6133: oled_colour = 16'b00000_000000_00000;
		6134: oled_colour = 16'b00000_000000_00000;
		6135: oled_colour = 16'b00000_000000_00000;
		6136: oled_colour = 16'b00000_000000_00000;
		6137: oled_colour = 16'b00000_000000_00000;
		6138: oled_colour = 16'b00000_000000_00000;
		6139: oled_colour = 16'b00000_000000_00000;
		6140: oled_colour = 16'b00000_000000_00000;
		6141: oled_colour = 16'b00000_000000_00000;
		6142: oled_colour = 16'b00000_000000_00000;
		6143: oled_colour = 16'b00000_000000_00000;
		default: oled_colour = 16'b00000_000000_00000; 
	endcase
end

endmodule