module Gui_Sp2(
    input [12:0] pixel_index, 
    output reg [15:0] oled_colour 
); 

always@(pixel_index) 
begin
	case(pixel_index)
		1675: oled_colour = 16'b01100_011110_11001; 
		1676: oled_colour = 16'b01101_100100_11011; 
		1677: oled_colour = 16'b10001_110001_11101; 
		1678: oled_colour = 16'b10100_110101_11101; 
		1765: oled_colour = 16'b10100_110001_11110; 
		1766: oled_colour = 16'b10110_110010_11110; 
		1767: oled_colour = 16'b11000_110111_11111; 
		1768: oled_colour = 16'b11011_111100_11111; 
		1769: oled_colour = 16'b11101_111110_11111; 
		1770: oled_colour = 16'b11101_111110_11111; 
		1771: oled_colour = 16'b11110_111100_11111; 
		1772: oled_colour = 16'b11110_111011_11111; 
		1773: oled_colour = 16'b11110_111100_11111; 
		1775: oled_colour = 16'b11110_111111_11111; 
		1776: oled_colour = 16'b11000_111011_11111; 
		1777: oled_colour = 16'b10000_110000_11111; 
		1778: oled_colour = 16'b01011_100110_11100; 
		1859: oled_colour = 16'b10100_101101_11010; 
		1860: oled_colour = 16'b11000_110110_11011; 
		1861: oled_colour = 16'b11110_111001_11001; 
		1862: oled_colour = 16'b11111_110111_11000; 
		1863: oled_colour = 16'b11111_111000_11000; 
		1864: oled_colour = 16'b11111_111010_11000; 
		1865: oled_colour = 16'b11111_111011_11010; 
		1866: oled_colour = 16'b11111_111011_11011; 
		1867: oled_colour = 16'b11111_111111_11101; 
		1868: oled_colour = 16'b11111_111111_11110; 
		1870: oled_colour = 16'b11111_111101_11111; 
		1871: oled_colour = 16'b11111_111011_11101; 
		1872: oled_colour = 16'b11111_111111_11101; 
		1873: oled_colour = 16'b11101_111001_11010; 
		1874: oled_colour = 16'b11100_110011_10011; 
		1875: oled_colour = 16'b11010_110001_01110; 
		1876: oled_colour = 16'b10100_101000_10011; 
		1965: oled_colour = 16'b11101_110010_10001; 
		1966: oled_colour = 16'b11101_110000_10001; 
		1967: oled_colour = 16'b11101_101110_01101; 
		1968: oled_colour = 16'b11101_110001_01100; 
		1969: oled_colour = 16'b11110_110110_00110; 
		1970: oled_colour = 16'b11110_110001_01000; 
		1971: oled_colour = 16'b11111_110011_01010; 
		1972: oled_colour = 16'b11110_111000_00111; 
		1973: oled_colour = 16'b11111_111010_01000; 
		2063: oled_colour = 16'b10101_100010_01100; 
		2064: oled_colour = 16'b10111_100011_01011; 
		2065: oled_colour = 16'b11110_110001_01011; 
		2066: oled_colour = 16'b11110_110111_00110; 
		2067: oled_colour = 16'b11101_101110_01101; 
		2068: oled_colour = 16'b11111_110110_01010; 
		2069: oled_colour = 16'b11111_110111_01010; 
		2070: oled_colour = 16'b01111_100101_10110; 
		2158: oled_colour = 16'b01001_011000_00101; 
		2159: oled_colour = 16'b10100_100000_01100; 
		2160: oled_colour = 16'b11100_101101_01111; 
		2161: oled_colour = 16'b11100_101110_01101; 
		2162: oled_colour = 16'b11101_101110_01100; 
		2163: oled_colour = 16'b11010_100111_01111; 
		2164: oled_colour = 16'b11010_101110_10100; 
		2165: oled_colour = 16'b11010_101110_10010; 
		2251: oled_colour = 16'b11001_101110_10001; 
		2252: oled_colour = 16'b11001_101110_10010; 
		2253: oled_colour = 16'b10100_100111_01111; 
		2254: oled_colour = 16'b11001_110010_10100; 
		2255: oled_colour = 16'b11010_101010_10001; 
		2256: oled_colour = 16'b11101_101101_10010; 
		2257: oled_colour = 16'b11010_101001_10000; 
		2258: oled_colour = 16'b11001_100010_01110; 
		2259: oled_colour = 16'b11101_101111_10010; 
		2260: oled_colour = 16'b11011_101110_10011; 
		2346: oled_colour = 16'b11101_101011_10000; 
		2347: oled_colour = 16'b11111_111111_11100; 
		2348: oled_colour = 16'b11111_111011_11100; 
		2349: oled_colour = 16'b11111_110101_11000; 
		2350: oled_colour = 16'b10111_110010_10100; 
		2351: oled_colour = 16'b10110_101001_01111; 
		2352: oled_colour = 16'b11010_100101_01111; 
		2353: oled_colour = 16'b11010_101010_10000; 
		2354: oled_colour = 16'b10110_011100_01010; 
		2355: oled_colour = 16'b11101_101101_10001; 
		2356: oled_colour = 16'b11010_101000_10000; 
		2441: oled_colour = 16'b11010_011011_01000; 
		2442: oled_colour = 16'b11001_100000_01110; 
		2443: oled_colour = 16'b11100_101100_10001; 
		2444: oled_colour = 16'b11111_110111_10110; 
		2445: oled_colour = 16'b11111_110111_10111; 
		2446: oled_colour = 16'b11010_101011_10001; 
		2447: oled_colour = 16'b10111_110100_10011; 
		2448: oled_colour = 16'b11001_100111_01110; 
		2449: oled_colour = 16'b11000_100010_01101; 
		2450: oled_colour = 16'b10110_100000_01100; 
		2451: oled_colour = 16'b10010_011011_01000; 
		2536: oled_colour = 16'b11100_101100_10001; 
		2537: oled_colour = 16'b11111_110001_10100; 
		2538: oled_colour = 16'b11011_100100_01110; 
		2539: oled_colour = 16'b11100_101001_10000; 
		2540: oled_colour = 16'b11001_100100_01101; 
		2541: oled_colour = 16'b11100_101010_01111; 
		2542: oled_colour = 16'b11111_110011_10100; 
		2543: oled_colour = 16'b10100_110111_10100; 
		2544: oled_colour = 16'b10100_110110_10011; 
		2545: oled_colour = 16'b11001_101101_10010; 
		2546: oled_colour = 16'b11000_100011_01101; 
		2547: oled_colour = 16'b10001_011111_01010; 
		2631: oled_colour = 16'b11100_101000_10000; 
		2632: oled_colour = 16'b11110_110000_10010; 
		2633: oled_colour = 16'b11110_110100_10110; 
		2634: oled_colour = 16'b11111_111000_11001; 
		2635: oled_colour = 16'b11001_100110_01110; 
		2636: oled_colour = 16'b10100_011001_01001; 
		2637: oled_colour = 16'b10101_011111_01011; 
		2638: oled_colour = 16'b10100_101000_01110; 
		2639: oled_colour = 16'b10000_101110_10001; 
		2640: oled_colour = 16'b10001_110101_10011; 
		2641: oled_colour = 16'b10100_110101_10101; 
		2642: oled_colour = 16'b10011_100110_01101; 
		2726: oled_colour = 16'b11111_110010_10011; 
		2727: oled_colour = 16'b11110_110000_10011; 
		2728: oled_colour = 16'b11100_101011_10001; 
		2729: oled_colour = 16'b10111_100000_01101; 
		2730: oled_colour = 16'b10001_011111_01010; 
		2731: oled_colour = 16'b00110_010101_00010; 
		2732: oled_colour = 16'b01101_011110_01000; 
		2733: oled_colour = 16'b01000_011010_00110; 
		2734: oled_colour = 16'b00110_011010_00110; 
		2735: oled_colour = 16'b01100_100011_01100; 
		2736: oled_colour = 16'b01100_100100_01100; 
		2737: oled_colour = 16'b01010_100000_01010; 
		2738: oled_colour = 16'b00110_011010_00111; 
		2819: oled_colour = 16'b10101_110101_11011; 
		2821: oled_colour = 16'b11100_110000_10010; 
		2822: oled_colour = 16'b11110_111010_10111; 
		2823: oled_colour = 16'b11110_111001_10110; 
		2824: oled_colour = 16'b11111_110011_10010; 
		2825: oled_colour = 16'b10110_100010_01010; 
		2826: oled_colour = 16'b00011_010000_00001; 
		2827: oled_colour = 16'b00001_010100_00001; 
		2828: oled_colour = 16'b00011_010111_00011; 
		2829: oled_colour = 16'b00100_010110_00010; 
		2830: oled_colour = 16'b00110_011000_00101; 
		2910: oled_colour = 16'b01010_100110_11100; 
		2911: oled_colour = 16'b10000_110010_11111; 
		2912: oled_colour = 16'b10110_111001_11110; 
		2913: oled_colour = 16'b11100_111101_11111; 
		2914: oled_colour = 16'b11101_111100_11110; 
		2915: oled_colour = 16'b11110_111110_11111; 
		2918: oled_colour = 16'b11111_111101_11110; 
		2919: oled_colour = 16'b11111_111101_11101; 
		2920: oled_colour = 16'b11110_111100_11001; 
		2921: oled_colour = 16'b11111_111011_10010; 
		2922: oled_colour = 16'b11100_110001_01001; 
		2923: oled_colour = 16'b10100_011110_00011; 
		2924: oled_colour = 16'b01101_010111_00100; 
		2925: oled_colour = 16'b10011_101001_10000; 
		3006: oled_colour = 16'b01001_100011_11010; 
		3007: oled_colour = 16'b01101_101100_11110; 
		3008: oled_colour = 16'b10100_110101_11111; 
		3009: oled_colour = 16'b11010_111011_11111; 
		3010: oled_colour = 16'b11101_111101_11111; 
		3011: oled_colour = 16'b11111_111101_11110; 
		3012: oled_colour = 16'b11111_111100_11110; 
		3013: oled_colour = 16'b11110_111100_11110; 
		3014: oled_colour = 16'b11111_111101_11111; 
		3015: oled_colour = 16'b11111_111101_11111; 
		3016: oled_colour = 16'b11110_111101_11111; 
		3017: oled_colour = 16'b11110_111101_11110; 
		3018: oled_colour = 16'b11101_111111_11011; 
		3019: oled_colour = 16'b11010_110110_10101; 
		3020: oled_colour = 16'b10000_100000_10001; 
		3021: oled_colour = 16'b01100_011111_01011; 
		3022: oled_colour = 16'b10010_011110_01001; 
		3105: oled_colour = 16'b10100_110011_11101; 
		3106: oled_colour = 16'b10111_111000_11111; 
		3107: oled_colour = 16'b11011_111100_11111; 
		3108: oled_colour = 16'b11111_111101_11111; 
		3109: oled_colour = 16'b11111_111101_11111; 
		3110: oled_colour = 16'b11111_111100_11110; 
		3111: oled_colour = 16'b11110_111100_11110; 
		3112: oled_colour = 16'b11111_111100_11110; 
		3113: oled_colour = 16'b11111_111101_11111; 
		3114: oled_colour = 16'b11101_111101_11111; 
		3115: oled_colour = 16'b10011_111000_11111; 
		3116: oled_colour = 16'b01100_101001_11101; 
		3117: oled_colour = 16'b00111_011000_00110; 
		3118: oled_colour = 16'b01111_011001_00111; 
		3119: oled_colour = 16'b10101_101001_01111; 
		3120: oled_colour = 16'b10110_110001_10010; 
		3121: oled_colour = 16'b11010_101011_10011; 
		3202: oled_colour = 16'b01111_101110_11101; 
		3203: oled_colour = 16'b10100_110101_11111; 
		3204: oled_colour = 16'b11011_111101_11111; 
		3205: oled_colour = 16'b11110_111111_11111; 
		3208: oled_colour = 16'b11110_111110_11111; 
		3209: oled_colour = 16'b11010_111100_11111; 
		3210: oled_colour = 16'b10011_110110_11111; 
		3211: oled_colour = 16'b01100_101011_11101; 
		3212: oled_colour = 16'b10011_101110_11010; 
		3213: oled_colour = 16'b01011_100000_01001; 
		3214: oled_colour = 16'b01011_010100_00100; 
		3215: oled_colour = 16'b10100_101101_10001; 
		3216: oled_colour = 16'b11111_111011_11001; 
		3217: oled_colour = 16'b11111_111000_10110; 
		3218: oled_colour = 16'b11111_101110_10001; 
		3219: oled_colour = 16'b11100_100110_01111; 
		3220: oled_colour = 16'b10110_011111_01011; 
		3304: oled_colour = 16'b11000_110001_11001; 
		3305: oled_colour = 16'b10010_101010_10111; 
		3306: oled_colour = 16'b10011_101001_11000; 
		3307: oled_colour = 16'b11010_101111_10110; 
		3308: oled_colour = 16'b11111_111011_11000; 
		3309: oled_colour = 16'b10010_101101_10000; 
		3310: oled_colour = 16'b01000_010110_00100; 
		3311: oled_colour = 16'b01110_101000_01111; 
		3312: oled_colour = 16'b10110_110111_10100; 
		3313: oled_colour = 16'b11010_111001_10100; 
		3314: oled_colour = 16'b11111_110001_10010; 
		3315: oled_colour = 16'b11100_110101_10011; 
		3316: oled_colour = 16'b11010_110111_10011; 
		3317: oled_colour = 16'b10111_110111_10011; 
		3401: oled_colour = 16'b11111_111001_11000; 
		3402: oled_colour = 16'b11100_110111_10111; 
		3403: oled_colour = 16'b11011_101110_01111; 
		3404: oled_colour = 16'b11111_110111_10101; 
		3405: oled_colour = 16'b10110_110011_10010; 
		3406: oled_colour = 16'b00100_010111_00100; 
		3407: oled_colour = 16'b01011_011100_01000; 
		3408: oled_colour = 16'b10101_101100_10010; 
		3409: oled_colour = 16'b01100_100011_01100; 
		3410: oled_colour = 16'b10000_101001_01101; 
		3411: oled_colour = 16'b01100_100110_01100; 
		3412: oled_colour = 16'b10011_110001_10010; 
		3413: oled_colour = 16'b11101_111110_10110; 
		3414: oled_colour = 16'b10000_100111_01100; 
		3497: oled_colour = 16'b10011_101111_10001; 
		3498: oled_colour = 16'b10010_110011_10100; 
		3499: oled_colour = 16'b10110_110110_10011; 
		3500: oled_colour = 16'b11110_111011_11010; 
		3501: oled_colour = 16'b11011_110110_10110; 
		3505: oled_colour = 16'b01000_010110_00100; 
		3506: oled_colour = 16'b10100_011100_01010; 
		3507: oled_colour = 16'b10101_101101_10001; 
		3508: oled_colour = 16'b11010_111110_10100; 
		3509: oled_colour = 16'b11000_110101_10010; 
		3510: oled_colour = 16'b01110_011011_01000; 
		3592: oled_colour = 16'b10011_011001_00111; 
		3593: oled_colour = 16'b01001_001111_00001; 
		3594: oled_colour = 16'b01100_100011_01011; 
		3595: oled_colour = 16'b11011_111100_11001; 
		3596: oled_colour = 16'b11111_111101_11111; 
		3597: oled_colour = 16'b11101_111111_11100; 
		3598: oled_colour = 16'b01101_100110_01101; 
		3601: oled_colour = 16'b01001_011101_00111; 
		3602: oled_colour = 16'b11000_110011_10100; 
		3603: oled_colour = 16'b11111_111000_11000; 
		3604: oled_colour = 16'b11110_111011_11000; 
		3605: oled_colour = 16'b10110_101111_10010; 
		3687: oled_colour = 16'b01101_011000_00110; 
		3688: oled_colour = 16'b11101_110101_11000; 
		3689: oled_colour = 16'b11010_101111_10001; 
		3690: oled_colour = 16'b10011_101001_01111; 
		3691: oled_colour = 16'b10110_101111_10010; 
		3692: oled_colour = 16'b11111_111110_11100; 
		3693: oled_colour = 16'b11001_111011_10111; 
		3697: oled_colour = 16'b01111_011101_01000; 
		3698: oled_colour = 16'b01010_100010_01010; 
		3699: oled_colour = 16'b10000_101000_01110; 
		3700: oled_colour = 16'b10011_100101_01111; 
		3782: oled_colour = 16'b10100_011110_01010; 
		3783: oled_colour = 16'b01010_011000_00100; 
		3784: oled_colour = 16'b11000_110000_10011; 
		3785: oled_colour = 16'b11111_111101_11100; 
		3786: oled_colour = 16'b11111_111011_11000; 
		3787: oled_colour = 16'b11011_110110_10011; 
		3788: oled_colour = 16'b10011_110000_10001; 
		3793: oled_colour = 16'b10011_011010_00110; 
		3794: oled_colour = 16'b10011_011101_01001; 
		3795: oled_colour = 16'b01110_011010_00111; 
		3876: oled_colour = 16'b10101_011101_01001; 
		3877: oled_colour = 16'b01011_001111_00001; 
		3878: oled_colour = 16'b10110_011110_01010; 
		3879: oled_colour = 16'b10010_011110_01000; 
		3880: oled_colour = 16'b01010_010111_00100; 
		3881: oled_colour = 16'b10110_101011_01111; 
		3888: oled_colour = 16'b01101_010001_00010; 
		3889: oled_colour = 16'b01110_010011_00010; 
		3890: oled_colour = 16'b10111_100000_01010; 
		3971: oled_colour = 16'b10110_011111_01100; 
		3972: oled_colour = 16'b01111_010100_00011; 
		3973: oled_colour = 16'b01111_010110_00100; 
		3974: oled_colour = 16'b10011_011001_00111; 
		3983: oled_colour = 16'b11001_100011_01101; 
		3984: oled_colour = 16'b01101_010010_00010; 
		3985: oled_colour = 16'b10011_011100_00111; 
		4068: oled_colour = 16'b01100_010001_00001; 
		4069: oled_colour = 16'b10000_011000_00101; 
		4070: oled_colour = 16'b10111_100010_01011; 
		4079: oled_colour = 16'b10110_011110_01010; 
		4080: oled_colour = 16'b01100_010000_00001; 
		4081: oled_colour = 16'b01111_010101_00011; 
		4082: oled_colour = 16'b10110_011110_01011; 
		4165: oled_colour = 16'b10111_100100_01011; 
		4166: oled_colour = 16'b11111_110111_10111; 
		4167: oled_colour = 16'b11010_100100_01110; 
		4178: oled_colour = 16'b11000_100000_01100; 
		4179: oled_colour = 16'b11101_101100_10001; 
		4180: oled_colour = 16'b11000_100010_01101; 
		default: oled_colour = 16'b00000_000000_00000; 
	endcase
end

endmodule