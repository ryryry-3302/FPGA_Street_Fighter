module Background(
    input [12:0] pixel_index, 
    output reg [15:0] oled_colour 
); 

always@(pixel_index) 
begin
	case(pixel_index)
		0: oled_colour = 16'b00010_000101_00111; 
		1: oled_colour = 16'b00010_000101_00111; 
		2: oled_colour = 16'b00010_000101_00111; 
		3: oled_colour = 16'b00010_000101_00111; 
		4: oled_colour = 16'b00010_000101_00111; 
		5: oled_colour = 16'b00010_000101_00111; 
		6: oled_colour = 16'b00010_000101_00111; 
		7: oled_colour = 16'b00010_000101_00111; 
		8: oled_colour = 16'b00010_000101_00111; 
		9: oled_colour = 16'b00010_000101_00111; 
		10: oled_colour = 16'b00010_000101_00111; 
		11: oled_colour = 16'b00010_000101_00111; 
		12: oled_colour = 16'b00010_000101_00111; 
		13: oled_colour = 16'b00010_000101_00111; 
		14: oled_colour = 16'b00010_000101_00111; 
		15: oled_colour = 16'b00010_000101_00111; 
		16: oled_colour = 16'b00010_000101_00111; 
		17: oled_colour = 16'b00010_000101_00111; 
		18: oled_colour = 16'b00010_000101_00111; 
		19: oled_colour = 16'b00010_000101_00111; 
		20: oled_colour = 16'b00010_000101_00111; 
		21: oled_colour = 16'b00010_000101_00111; 
		22: oled_colour = 16'b00010_000101_00111; 
		23: oled_colour = 16'b00010_000101_00111; 
		24: oled_colour = 16'b00010_000101_00111; 
		25: oled_colour = 16'b00010_000101_00111; 
		26: oled_colour = 16'b00010_000101_00111; 
		27: oled_colour = 16'b00010_000101_00111; 
		28: oled_colour = 16'b00010_000101_00111; 
		29: oled_colour = 16'b00010_000101_00111; 
		30: oled_colour = 16'b00010_000101_00111; 
		31: oled_colour = 16'b00010_000101_00111; 
		32: oled_colour = 16'b00010_000101_00111; 
		33: oled_colour = 16'b00010_000101_00111; 
		34: oled_colour = 16'b00010_000101_00111; 
		35: oled_colour = 16'b00010_000101_00111; 
		36: oled_colour = 16'b00010_000101_00111; 
		37: oled_colour = 16'b00010_000101_00111; 
		38: oled_colour = 16'b00010_000101_00111; 
		39: oled_colour = 16'b00010_000101_00111; 
		40: oled_colour = 16'b00010_000101_00111; 
		41: oled_colour = 16'b00010_000101_00111; 
		42: oled_colour = 16'b00010_000101_00111; 
		43: oled_colour = 16'b00010_000101_00111; 
		44: oled_colour = 16'b00010_000101_00111; 
		45: oled_colour = 16'b00010_000101_00111; 
		46: oled_colour = 16'b00010_000101_00111; 
		47: oled_colour = 16'b00010_000101_00111; 
		48: oled_colour = 16'b00010_000101_00111; 
		49: oled_colour = 16'b00010_000101_00111; 
		50: oled_colour = 16'b00010_000101_00111; 
		51: oled_colour = 16'b00010_000101_00111; 
		52: oled_colour = 16'b00010_000101_00111; 
		53: oled_colour = 16'b00010_000101_00111; 
		54: oled_colour = 16'b00010_000101_00111; 
		55: oled_colour = 16'b00010_000101_00111; 
		56: oled_colour = 16'b00010_000101_00111; 
		57: oled_colour = 16'b00010_000101_00111; 
		58: oled_colour = 16'b00010_000101_00111; 
		59: oled_colour = 16'b00010_000101_00111; 
		60: oled_colour = 16'b00010_000101_00111; 
		61: oled_colour = 16'b00010_000101_00111; 
		62: oled_colour = 16'b00010_000101_00111; 
		63: oled_colour = 16'b00010_000101_00111; 
		64: oled_colour = 16'b00010_000101_00111; 
		65: oled_colour = 16'b00010_000101_00111; 
		66: oled_colour = 16'b00010_000101_00111; 
		67: oled_colour = 16'b00010_000101_00111; 
		68: oled_colour = 16'b00010_000101_00111; 
		69: oled_colour = 16'b00010_000101_00111; 
		70: oled_colour = 16'b00010_000101_00111; 
		71: oled_colour = 16'b00010_000101_00111; 
		72: oled_colour = 16'b00010_000101_00111; 
		73: oled_colour = 16'b00010_000101_00111; 
		74: oled_colour = 16'b00010_000101_00111; 
		75: oled_colour = 16'b00010_000101_00111; 
		76: oled_colour = 16'b00010_000101_00111; 
		77: oled_colour = 16'b00010_000101_00111; 
		78: oled_colour = 16'b00010_000101_00111; 
		79: oled_colour = 16'b00010_000101_00111; 
		80: oled_colour = 16'b00010_000101_00111; 
		81: oled_colour = 16'b00010_000101_00111; 
		82: oled_colour = 16'b00010_000101_00111; 
		83: oled_colour = 16'b00010_000101_00111; 
		84: oled_colour = 16'b00010_000101_00111; 
		85: oled_colour = 16'b00010_000101_00111; 
		86: oled_colour = 16'b00010_000101_00111; 
		87: oled_colour = 16'b00010_000101_00111; 
		88: oled_colour = 16'b00010_000101_00111; 
		89: oled_colour = 16'b00010_000101_00111; 
		90: oled_colour = 16'b00010_000101_00111; 
		91: oled_colour = 16'b00010_000101_00111; 
		92: oled_colour = 16'b00010_000101_00111; 
		93: oled_colour = 16'b00010_000101_00111; 
		94: oled_colour = 16'b00010_000101_00111; 
		95: oled_colour = 16'b00010_000101_00111; 
		96: oled_colour = 16'b00010_000101_00111; 
		97: oled_colour = 16'b00010_000101_00111; 
		98: oled_colour = 16'b00010_000101_00111; 
		99: oled_colour = 16'b00010_000101_00111; 
		100: oled_colour = 16'b00010_000101_00111; 
		101: oled_colour = 16'b00010_000101_00111; 
		102: oled_colour = 16'b00010_000101_00111; 
		103: oled_colour = 16'b00010_000101_00111; 
		104: oled_colour = 16'b00010_000101_00111; 
		105: oled_colour = 16'b00010_000101_00111; 
		106: oled_colour = 16'b00010_000101_00111; 
		107: oled_colour = 16'b00010_000101_00111; 
		108: oled_colour = 16'b00010_000101_00111; 
		109: oled_colour = 16'b00010_000101_00111; 
		110: oled_colour = 16'b00010_000101_00111; 
		111: oled_colour = 16'b00010_000101_00111; 
		112: oled_colour = 16'b00010_000101_00111; 
		113: oled_colour = 16'b00010_000101_00111; 
		114: oled_colour = 16'b00010_000101_00111; 
		115: oled_colour = 16'b00010_000101_00111; 
		116: oled_colour = 16'b00010_000101_00111; 
		117: oled_colour = 16'b00010_000101_00111; 
		118: oled_colour = 16'b00010_000101_00111; 
		119: oled_colour = 16'b00010_000101_00111; 
		120: oled_colour = 16'b00010_000101_00111; 
		121: oled_colour = 16'b00010_000101_00111; 
		122: oled_colour = 16'b00010_000101_00111; 
		123: oled_colour = 16'b00010_000101_00111; 
		124: oled_colour = 16'b00010_000101_00111; 
		125: oled_colour = 16'b00010_000101_00111; 
		126: oled_colour = 16'b00010_000101_00111; 
		127: oled_colour = 16'b00010_000101_00111; 
		128: oled_colour = 16'b00010_000101_00111; 
		129: oled_colour = 16'b00010_000101_00111; 
		130: oled_colour = 16'b00010_000101_00111; 
		131: oled_colour = 16'b00010_000101_00111; 
		132: oled_colour = 16'b00010_000101_00111; 
		133: oled_colour = 16'b00010_000101_00111; 
		134: oled_colour = 16'b00010_000101_00111; 
		135: oled_colour = 16'b00010_000101_00111; 
		136: oled_colour = 16'b00010_000101_00111; 
		137: oled_colour = 16'b00010_000101_00111; 
		138: oled_colour = 16'b00010_000101_00111; 
		139: oled_colour = 16'b00010_000101_00111; 
		140: oled_colour = 16'b00010_000101_00111; 
		141: oled_colour = 16'b00010_000101_00111; 
		142: oled_colour = 16'b00010_000101_00111; 
		143: oled_colour = 16'b00010_000101_00111; 
		144: oled_colour = 16'b00010_000101_00111; 
		145: oled_colour = 16'b00010_000101_00111; 
		146: oled_colour = 16'b00010_000101_00111; 
		147: oled_colour = 16'b00010_000101_00111; 
		148: oled_colour = 16'b00010_000101_00111; 
		149: oled_colour = 16'b00010_000101_00111; 
		150: oled_colour = 16'b00010_000101_00111; 
		151: oled_colour = 16'b00010_000101_00111; 
		152: oled_colour = 16'b00010_000101_00111; 
		153: oled_colour = 16'b00010_000101_00111; 
		154: oled_colour = 16'b00010_000101_00111; 
		155: oled_colour = 16'b00010_000101_00111; 
		156: oled_colour = 16'b00010_000101_00111; 
		157: oled_colour = 16'b00010_000101_00111; 
		158: oled_colour = 16'b00010_000101_00111; 
		159: oled_colour = 16'b00010_000101_00111; 
		160: oled_colour = 16'b00010_000101_00111; 
		161: oled_colour = 16'b00010_000101_00111; 
		162: oled_colour = 16'b00010_000101_00111; 
		163: oled_colour = 16'b00010_000101_00111; 
		164: oled_colour = 16'b00010_000101_00111; 
		165: oled_colour = 16'b00010_000101_00111; 
		166: oled_colour = 16'b00010_000101_00111; 
		167: oled_colour = 16'b00010_000101_00111; 
		168: oled_colour = 16'b00010_000101_00111; 
		169: oled_colour = 16'b00010_000101_00111; 
		170: oled_colour = 16'b00010_000101_00111; 
		171: oled_colour = 16'b00010_000101_00111; 
		172: oled_colour = 16'b00010_000101_00111; 
		173: oled_colour = 16'b00010_000101_00111; 
		174: oled_colour = 16'b00010_000101_00111; 
		175: oled_colour = 16'b00010_000101_00111; 
		176: oled_colour = 16'b00010_000101_00111; 
		177: oled_colour = 16'b00010_000101_00111; 
		178: oled_colour = 16'b00010_000101_00111; 
		179: oled_colour = 16'b00010_000101_00111; 
		180: oled_colour = 16'b00010_000101_00111; 
		181: oled_colour = 16'b00010_000101_00111; 
		182: oled_colour = 16'b00011_000101_00111; 
		183: oled_colour = 16'b00011_000101_00111; 
		184: oled_colour = 16'b00010_000101_00111; 
		185: oled_colour = 16'b00010_000101_00111; 
		186: oled_colour = 16'b00010_000101_00111; 
		187: oled_colour = 16'b00010_000101_00111; 
		188: oled_colour = 16'b00010_000101_00111; 
		189: oled_colour = 16'b00010_000101_00111; 
		190: oled_colour = 16'b00010_000101_00111; 
		191: oled_colour = 16'b00010_000101_00111; 
		192: oled_colour = 16'b00010_000101_00111; 
		193: oled_colour = 16'b00010_000101_00111; 
		194: oled_colour = 16'b00010_000101_00111; 
		195: oled_colour = 16'b00010_000101_00111; 
		196: oled_colour = 16'b00010_000101_00111; 
		197: oled_colour = 16'b00010_000101_00111; 
		198: oled_colour = 16'b00010_000101_00111; 
		199: oled_colour = 16'b00010_000101_00111; 
		200: oled_colour = 16'b00010_000101_00111; 
		201: oled_colour = 16'b00011_000101_00111; 
		202: oled_colour = 16'b00011_000101_00111; 
		203: oled_colour = 16'b00011_000101_00111; 
		204: oled_colour = 16'b00010_000101_00111; 
		205: oled_colour = 16'b00010_000101_00111; 
		206: oled_colour = 16'b00010_000101_00111; 
		207: oled_colour = 16'b00010_000101_00111; 
		208: oled_colour = 16'b00010_000101_00111; 
		209: oled_colour = 16'b00010_000101_00111; 
		210: oled_colour = 16'b00010_000101_00111; 
		211: oled_colour = 16'b00010_000101_00111; 
		212: oled_colour = 16'b00010_000101_00111; 
		213: oled_colour = 16'b00010_000101_00111; 
		214: oled_colour = 16'b00010_000101_00111; 
		215: oled_colour = 16'b00010_000101_00111; 
		216: oled_colour = 16'b00010_000101_00111; 
		217: oled_colour = 16'b00010_000101_00111; 
		218: oled_colour = 16'b00010_000101_00111; 
		219: oled_colour = 16'b00010_000101_00111; 
		220: oled_colour = 16'b00010_000101_00111; 
		221: oled_colour = 16'b00010_000101_00111; 
		222: oled_colour = 16'b00010_000101_00111; 
		223: oled_colour = 16'b00010_000101_00111; 
		224: oled_colour = 16'b00010_000101_00111; 
		225: oled_colour = 16'b00010_000101_00111; 
		226: oled_colour = 16'b00010_000101_00111; 
		227: oled_colour = 16'b00010_000101_00111; 
		228: oled_colour = 16'b00010_000101_00111; 
		229: oled_colour = 16'b00010_000101_00111; 
		230: oled_colour = 16'b00010_000101_00111; 
		231: oled_colour = 16'b00010_000101_00111; 
		232: oled_colour = 16'b00010_000101_00111; 
		233: oled_colour = 16'b00010_000101_00111; 
		234: oled_colour = 16'b00010_000101_00111; 
		235: oled_colour = 16'b00010_000101_00111; 
		236: oled_colour = 16'b00010_000101_00111; 
		237: oled_colour = 16'b00010_000101_00111; 
		238: oled_colour = 16'b00010_000101_00111; 
		239: oled_colour = 16'b00010_000101_00111; 
		240: oled_colour = 16'b00010_000101_00111; 
		241: oled_colour = 16'b00010_000101_00111; 
		242: oled_colour = 16'b00010_000101_00111; 
		243: oled_colour = 16'b00010_000101_00111; 
		244: oled_colour = 16'b00010_000101_00111; 
		245: oled_colour = 16'b00010_000101_00111; 
		246: oled_colour = 16'b00010_000101_00111; 
		247: oled_colour = 16'b00010_000101_00111; 
		248: oled_colour = 16'b00010_000101_00111; 
		249: oled_colour = 16'b00010_000101_00111; 
		250: oled_colour = 16'b00010_000101_00111; 
		251: oled_colour = 16'b00010_000101_00111; 
		252: oled_colour = 16'b00010_000101_00111; 
		253: oled_colour = 16'b00010_000101_00111; 
		254: oled_colour = 16'b00010_000101_00111; 
		255: oled_colour = 16'b00010_000101_00111; 
		256: oled_colour = 16'b00010_000101_00111; 
		257: oled_colour = 16'b00010_000101_00111; 
		258: oled_colour = 16'b00010_000101_00111; 
		259: oled_colour = 16'b00010_000101_00111; 
		260: oled_colour = 16'b00010_000101_00111; 
		261: oled_colour = 16'b00010_000101_00111; 
		262: oled_colour = 16'b00010_000101_00111; 
		263: oled_colour = 16'b00010_000101_00111; 
		264: oled_colour = 16'b00010_000101_00111; 
		265: oled_colour = 16'b00010_000101_00111; 
		266: oled_colour = 16'b00010_000101_00111; 
		267: oled_colour = 16'b00010_000101_00111; 
		268: oled_colour = 16'b00010_000101_00111; 
		269: oled_colour = 16'b00010_000101_00111; 
		270: oled_colour = 16'b00010_000101_00111; 
		271: oled_colour = 16'b00010_000101_00111; 
		272: oled_colour = 16'b00010_000101_00111; 
		273: oled_colour = 16'b00010_000101_00111; 
		274: oled_colour = 16'b00010_000101_00111; 
		275: oled_colour = 16'b00010_000101_00111; 
		276: oled_colour = 16'b00010_000101_00111; 
		277: oled_colour = 16'b00011_000111_00111; 
		278: oled_colour = 16'b00010_000100_00110; 
		279: oled_colour = 16'b00010_000101_00111; 
		280: oled_colour = 16'b00011_000110_00111; 
		281: oled_colour = 16'b00011_000101_00111; 
		282: oled_colour = 16'b00010_000101_00111; 
		283: oled_colour = 16'b00010_000101_00111; 
		284: oled_colour = 16'b00010_000101_00111; 
		285: oled_colour = 16'b00010_000101_00111; 
		286: oled_colour = 16'b00010_000101_00111; 
		287: oled_colour = 16'b00010_000101_00111; 
		288: oled_colour = 16'b00011_000101_00110; 
		289: oled_colour = 16'b00011_000101_00111; 
		290: oled_colour = 16'b00011_000101_00111; 
		291: oled_colour = 16'b00011_000101_00111; 
		292: oled_colour = 16'b00011_000101_00111; 
		293: oled_colour = 16'b00011_000101_00111; 
		294: oled_colour = 16'b00010_000101_00111; 
		295: oled_colour = 16'b00011_000101_00111; 
		296: oled_colour = 16'b00011_000101_00111; 
		297: oled_colour = 16'b00011_000100_00111; 
		298: oled_colour = 16'b00010_000100_00111; 
		299: oled_colour = 16'b00010_000100_00111; 
		300: oled_colour = 16'b00010_000100_00111; 
		301: oled_colour = 16'b00010_000101_00110; 
		302: oled_colour = 16'b00010_000101_00110; 
		303: oled_colour = 16'b00010_000101_00110; 
		304: oled_colour = 16'b00011_000101_00111; 
		305: oled_colour = 16'b00011_000101_00111; 
		306: oled_colour = 16'b00010_000101_00110; 
		307: oled_colour = 16'b00010_000101_00111; 
		308: oled_colour = 16'b00010_000101_00111; 
		309: oled_colour = 16'b00010_000101_00111; 
		310: oled_colour = 16'b00010_000101_00111; 
		311: oled_colour = 16'b00010_000101_00111; 
		312: oled_colour = 16'b00010_000101_00111; 
		313: oled_colour = 16'b00010_000101_00111; 
		314: oled_colour = 16'b00010_000101_00111; 
		315: oled_colour = 16'b00010_000101_00111; 
		316: oled_colour = 16'b00010_000101_00111; 
		317: oled_colour = 16'b00010_000101_00111; 
		318: oled_colour = 16'b00010_000101_00111; 
		319: oled_colour = 16'b00010_000101_00111; 
		320: oled_colour = 16'b00010_000101_00111; 
		321: oled_colour = 16'b00010_000101_00111; 
		322: oled_colour = 16'b00010_000101_00111; 
		323: oled_colour = 16'b00010_000101_00111; 
		324: oled_colour = 16'b00010_000101_00111; 
		325: oled_colour = 16'b00010_000101_00111; 
		326: oled_colour = 16'b00010_000101_00111; 
		327: oled_colour = 16'b00010_000101_00111; 
		328: oled_colour = 16'b00010_000101_00111; 
		329: oled_colour = 16'b00010_000101_00111; 
		330: oled_colour = 16'b00010_000101_00111; 
		331: oled_colour = 16'b00010_000101_00111; 
		332: oled_colour = 16'b00010_000101_00111; 
		333: oled_colour = 16'b00010_000101_00111; 
		334: oled_colour = 16'b00010_000101_00111; 
		335: oled_colour = 16'b00010_000101_00111; 
		336: oled_colour = 16'b00010_000101_00111; 
		337: oled_colour = 16'b00010_000101_00111; 
		338: oled_colour = 16'b00010_000101_00111; 
		339: oled_colour = 16'b00010_000101_00111; 
		340: oled_colour = 16'b00010_000101_00111; 
		341: oled_colour = 16'b00010_000101_00111; 
		342: oled_colour = 16'b00010_000101_00111; 
		343: oled_colour = 16'b00010_000101_00111; 
		344: oled_colour = 16'b00010_000101_00111; 
		345: oled_colour = 16'b00010_000101_00111; 
		346: oled_colour = 16'b00010_000101_00111; 
		347: oled_colour = 16'b00010_000101_00111; 
		348: oled_colour = 16'b00010_000101_00111; 
		349: oled_colour = 16'b00010_000101_00111; 
		350: oled_colour = 16'b00010_000101_00111; 
		351: oled_colour = 16'b00010_000101_00111; 
		352: oled_colour = 16'b00010_000101_00111; 
		353: oled_colour = 16'b00011_000101_00111; 
		354: oled_colour = 16'b00011_000101_00111; 
		355: oled_colour = 16'b00011_000101_00111; 
		356: oled_colour = 16'b00011_000101_00111; 
		357: oled_colour = 16'b00011_000101_00111; 
		358: oled_colour = 16'b00011_000101_00111; 
		359: oled_colour = 16'b00011_000101_00111; 
		360: oled_colour = 16'b00011_000101_00111; 
		361: oled_colour = 16'b00011_000101_00111; 
		362: oled_colour = 16'b00011_000101_00111; 
		363: oled_colour = 16'b00011_000101_00110; 
		364: oled_colour = 16'b00010_000101_00110; 
		365: oled_colour = 16'b00011_000101_00111; 
		366: oled_colour = 16'b00011_000101_00111; 
		367: oled_colour = 16'b00011_000101_00110; 
		368: oled_colour = 16'b00011_000101_00111; 
		369: oled_colour = 16'b00011_000101_00110; 
		370: oled_colour = 16'b00011_000101_00111; 
		371: oled_colour = 16'b00010_000100_00110; 
		372: oled_colour = 16'b00101_001010_01001; 
		373: oled_colour = 16'b01001_010100_01100; 
		374: oled_colour = 16'b01010_010100_01100; 
		375: oled_colour = 16'b00010_000100_00111; 
		376: oled_colour = 16'b00010_000011_00110; 
		377: oled_colour = 16'b00011_000101_00111; 
		378: oled_colour = 16'b00011_000101_00111; 
		379: oled_colour = 16'b00011_000101_00111; 
		380: oled_colour = 16'b00010_000101_00111; 
		381: oled_colour = 16'b00010_000101_00111; 
		382: oled_colour = 16'b00010_000101_00110; 
		383: oled_colour = 16'b00010_000101_00110; 
		384: oled_colour = 16'b00010_000101_01000; 
		385: oled_colour = 16'b00010_000101_01000; 
		386: oled_colour = 16'b00010_000101_01001; 
		387: oled_colour = 16'b00010_000101_01001; 
		388: oled_colour = 16'b00010_000110_01001; 
		389: oled_colour = 16'b00010_000111_01010; 
		390: oled_colour = 16'b00010_000111_01010; 
		391: oled_colour = 16'b00010_000111_01010; 
		392: oled_colour = 16'b00010_000111_01011; 
		393: oled_colour = 16'b00010_001000_01011; 
		394: oled_colour = 16'b00011_001000_01011; 
		395: oled_colour = 16'b00011_001001_01011; 
		396: oled_colour = 16'b00011_001001_01010; 
		397: oled_colour = 16'b00011_001000_01001; 
		398: oled_colour = 16'b00011_000110_01000; 
		399: oled_colour = 16'b00010_000110_01000; 
		400: oled_colour = 16'b00010_000110_01001; 
		401: oled_colour = 16'b00010_000101_01000; 
		402: oled_colour = 16'b00010_000101_01000; 
		403: oled_colour = 16'b00010_000101_01000; 
		404: oled_colour = 16'b00010_000101_00111; 
		405: oled_colour = 16'b00010_000101_00111; 
		406: oled_colour = 16'b00010_000101_00111; 
		407: oled_colour = 16'b00010_000101_00111; 
		408: oled_colour = 16'b00010_000101_00111; 
		409: oled_colour = 16'b00010_000101_00111; 
		410: oled_colour = 16'b00010_000101_00111; 
		411: oled_colour = 16'b00010_000101_00111; 
		412: oled_colour = 16'b00011_000101_00111; 
		413: oled_colour = 16'b00011_000110_00110; 
		414: oled_colour = 16'b00011_000101_00111; 
		415: oled_colour = 16'b00011_000101_00111; 
		416: oled_colour = 16'b00010_000101_00111; 
		417: oled_colour = 16'b00010_000101_00111; 
		418: oled_colour = 16'b00010_000101_00111; 
		419: oled_colour = 16'b00010_000101_00111; 
		420: oled_colour = 16'b00010_000101_00111; 
		421: oled_colour = 16'b00010_000101_00111; 
		422: oled_colour = 16'b00010_000101_00111; 
		423: oled_colour = 16'b00010_000101_00111; 
		424: oled_colour = 16'b00010_000101_00111; 
		425: oled_colour = 16'b00010_000101_00111; 
		426: oled_colour = 16'b00010_000101_00111; 
		427: oled_colour = 16'b00010_000101_00111; 
		428: oled_colour = 16'b00010_000101_00111; 
		429: oled_colour = 16'b00010_000101_00111; 
		430: oled_colour = 16'b00010_000101_00111; 
		431: oled_colour = 16'b00010_000101_00111; 
		432: oled_colour = 16'b00010_000101_00111; 
		433: oled_colour = 16'b00010_000101_00111; 
		434: oled_colour = 16'b00010_000101_00111; 
		435: oled_colour = 16'b00010_000101_00111; 
		436: oled_colour = 16'b00010_000101_00111; 
		437: oled_colour = 16'b00010_000101_00111; 
		438: oled_colour = 16'b00010_000101_00111; 
		439: oled_colour = 16'b00010_000101_00111; 
		440: oled_colour = 16'b00010_000101_00111; 
		441: oled_colour = 16'b00010_000101_00111; 
		442: oled_colour = 16'b00010_000101_00111; 
		443: oled_colour = 16'b00010_000101_00111; 
		444: oled_colour = 16'b00010_000101_00111; 
		445: oled_colour = 16'b00010_000101_00111; 
		446: oled_colour = 16'b00010_000101_00111; 
		447: oled_colour = 16'b00010_000101_00111; 
		448: oled_colour = 16'b00010_000101_01000; 
		449: oled_colour = 16'b00010_000100_01000; 
		450: oled_colour = 16'b00010_000100_01000; 
		451: oled_colour = 16'b00010_000100_00111; 
		452: oled_colour = 16'b00010_000100_00111; 
		453: oled_colour = 16'b00010_000100_00111; 
		454: oled_colour = 16'b00010_000100_01000; 
		455: oled_colour = 16'b00010_000100_01001; 
		456: oled_colour = 16'b00010_000100_01001; 
		457: oled_colour = 16'b00010_000101_01000; 
		458: oled_colour = 16'b00010_000101_01001; 
		459: oled_colour = 16'b00010_000101_01001; 
		460: oled_colour = 16'b00010_000101_01001; 
		461: oled_colour = 16'b00010_000101_01001; 
		462: oled_colour = 16'b00010_000101_01000; 
		463: oled_colour = 16'b00010_000101_01000; 
		464: oled_colour = 16'b00010_000101_01000; 
		465: oled_colour = 16'b00010_000101_01000; 
		466: oled_colour = 16'b00010_000101_01001; 
		467: oled_colour = 16'b00001_000011_01000; 
		468: oled_colour = 16'b00110_001100_01011; 
		469: oled_colour = 16'b00111_010001_01010; 
		470: oled_colour = 16'b10001_100101_10000; 
		471: oled_colour = 16'b10001_100010_10000; 
		472: oled_colour = 16'b00110_001100_01001; 
		473: oled_colour = 16'b00010_000101_01001; 
		474: oled_colour = 16'b00010_000110_01010; 
		475: oled_colour = 16'b00010_000110_01010; 
		476: oled_colour = 16'b00010_000110_01010; 
		477: oled_colour = 16'b00010_000110_01010; 
		478: oled_colour = 16'b00010_000110_01010; 
		479: oled_colour = 16'b00010_000110_01010; 
		480: oled_colour = 16'b00101_010001_01110; 
		481: oled_colour = 16'b00110_010001_01110; 
		482: oled_colour = 16'b00110_010010_01111; 
		483: oled_colour = 16'b00111_010011_10000; 
		484: oled_colour = 16'b00111_010100_10000; 
		485: oled_colour = 16'b00111_010101_10000; 
		486: oled_colour = 16'b00111_010101_10000; 
		487: oled_colour = 16'b00111_010101_10000; 
		488: oled_colour = 16'b00111_010101_10000; 
		489: oled_colour = 16'b01000_010111_10000; 
		490: oled_colour = 16'b01000_010111_10001; 
		491: oled_colour = 16'b01001_011000_10010; 
		492: oled_colour = 16'b01001_011000_10010; 
		493: oled_colour = 16'b01001_011000_10001; 
		494: oled_colour = 16'b01001_010111_10001; 
		495: oled_colour = 16'b01000_010101_10001; 
		496: oled_colour = 16'b00111_010100_10000; 
		497: oled_colour = 16'b00110_010001_01111; 
		498: oled_colour = 16'b00100_001110_01110; 
		499: oled_colour = 16'b00011_001010_01100; 
		500: oled_colour = 16'b00011_000110_01001; 
		501: oled_colour = 16'b00010_000101_00111; 
		502: oled_colour = 16'b00010_000101_00110; 
		503: oled_colour = 16'b00010_000100_00110; 
		504: oled_colour = 16'b00010_000101_00110; 
		505: oled_colour = 16'b00011_000101_00111; 
		506: oled_colour = 16'b00010_000101_00111; 
		507: oled_colour = 16'b00011_000101_00111; 
		508: oled_colour = 16'b00010_000100_00111; 
		509: oled_colour = 16'b00001_000011_01001; 
		510: oled_colour = 16'b00001_000100_01010; 
		511: oled_colour = 16'b00010_000111_01011; 
		512: oled_colour = 16'b00010_000110_01010; 
		513: oled_colour = 16'b00010_000101_01000; 
		514: oled_colour = 16'b00010_000101_00111; 
		515: oled_colour = 16'b00010_000101_00111; 
		516: oled_colour = 16'b00010_000101_00111; 
		517: oled_colour = 16'b00010_000101_00111; 
		518: oled_colour = 16'b00010_000101_00111; 
		519: oled_colour = 16'b00010_000101_00111; 
		520: oled_colour = 16'b00010_000101_00111; 
		521: oled_colour = 16'b00010_000101_00111; 
		522: oled_colour = 16'b00010_000101_00111; 
		523: oled_colour = 16'b00010_000101_00111; 
		524: oled_colour = 16'b00010_000101_00111; 
		525: oled_colour = 16'b00010_000101_00111; 
		526: oled_colour = 16'b00010_000101_00111; 
		527: oled_colour = 16'b00010_000101_00111; 
		528: oled_colour = 16'b00010_000101_00111; 
		529: oled_colour = 16'b00010_000101_00111; 
		530: oled_colour = 16'b00010_000101_00111; 
		531: oled_colour = 16'b00010_000101_00111; 
		532: oled_colour = 16'b00010_000101_00111; 
		533: oled_colour = 16'b00010_000101_00111; 
		534: oled_colour = 16'b00010_000101_00111; 
		535: oled_colour = 16'b00010_000101_00111; 
		536: oled_colour = 16'b00010_000101_00111; 
		537: oled_colour = 16'b00010_000101_00111; 
		538: oled_colour = 16'b00010_000101_00111; 
		539: oled_colour = 16'b00010_000101_00111; 
		540: oled_colour = 16'b00010_000101_00111; 
		541: oled_colour = 16'b00011_000101_01000; 
		542: oled_colour = 16'b00011_000101_01001; 
		543: oled_colour = 16'b00010_000101_01010; 
		544: oled_colour = 16'b00011_001000_01100; 
		545: oled_colour = 16'b00100_001011_01101; 
		546: oled_colour = 16'b00100_001100_01101; 
		547: oled_colour = 16'b00100_001100_01101; 
		548: oled_colour = 16'b00100_001101_01101; 
		549: oled_colour = 16'b00100_001101_01101; 
		550: oled_colour = 16'b00100_001101_01101; 
		551: oled_colour = 16'b00100_001101_01101; 
		552: oled_colour = 16'b00100_001110_01110; 
		553: oled_colour = 16'b00101_001111_01110; 
		554: oled_colour = 16'b00101_001111_01110; 
		555: oled_colour = 16'b00101_001111_01110; 
		556: oled_colour = 16'b00100_001111_01110; 
		557: oled_colour = 16'b00100_001101_01101; 
		558: oled_colour = 16'b00100_001101_01101; 
		559: oled_colour = 16'b00101_001111_01110; 
		560: oled_colour = 16'b00101_001111_01110; 
		561: oled_colour = 16'b00101_001111_01110; 
		562: oled_colour = 16'b00101_001111_01110; 
		563: oled_colour = 16'b00100_001110_01110; 
		564: oled_colour = 16'b00111_010010_01110; 
		565: oled_colour = 16'b00111_010000_01011; 
		566: oled_colour = 16'b00110_010000_01010; 
		567: oled_colour = 16'b01101_011101_01110; 
		568: oled_colour = 16'b10101_101011_10001; 
		569: oled_colour = 16'b01110_100000_01111; 
		570: oled_colour = 16'b01000_010110_01111; 
		571: oled_colour = 16'b01001_011000_01111; 
		572: oled_colour = 16'b00110_010010_01110; 
		573: oled_colour = 16'b00110_010011_01111; 
		574: oled_colour = 16'b00101_010000_01110; 
		575: oled_colour = 16'b00100_001111_01110; 
		576: oled_colour = 16'b00111_010101_01111; 
		577: oled_colour = 16'b01000_010111_10000; 
		578: oled_colour = 16'b01000_010111_10000; 
		579: oled_colour = 16'b00111_010101_10000; 
		580: oled_colour = 16'b00110_010010_01111; 
		581: oled_colour = 16'b00101_010001_01110; 
		582: oled_colour = 16'b00101_001110_01101; 
		583: oled_colour = 16'b00101_001101_01110; 
		584: oled_colour = 16'b00101_001100_01101; 
		585: oled_colour = 16'b00101_001100_01101; 
		586: oled_colour = 16'b00101_001100_01100; 
		587: oled_colour = 16'b00100_001011_01011; 
		588: oled_colour = 16'b00100_001011_01100; 
		589: oled_colour = 16'b00100_001010_01100; 
		590: oled_colour = 16'b00100_001010_01011; 
		591: oled_colour = 16'b00011_001011_01011; 
		592: oled_colour = 16'b00100_001010_01011; 
		593: oled_colour = 16'b00011_001001_01011; 
		594: oled_colour = 16'b00011_001000_01010; 
		595: oled_colour = 16'b00010_000111_01010; 
		596: oled_colour = 16'b00010_000110_01010; 
		597: oled_colour = 16'b00011_000111_01010; 
		598: oled_colour = 16'b00011_001001_01010; 
		599: oled_colour = 16'b00011_001001_01010; 
		600: oled_colour = 16'b00011_001000_01010; 
		601: oled_colour = 16'b00011_000110_01001; 
		602: oled_colour = 16'b00011_000110_01000; 
		603: oled_colour = 16'b00001_000100_01001; 
		604: oled_colour = 16'b00100_001100_01101; 
		605: oled_colour = 16'b01101_011011_01110; 
		606: oled_colour = 16'b10100_100111_01101; 
		607: oled_colour = 16'b10010_100101_01111; 
		608: oled_colour = 16'b00110_010011_01111; 
		609: oled_colour = 16'b00010_001000_01100; 
		610: oled_colour = 16'b00011_000110_01010; 
		611: oled_colour = 16'b00011_000101_01000; 
		612: oled_colour = 16'b00010_000101_00111; 
		613: oled_colour = 16'b00010_000101_00111; 
		614: oled_colour = 16'b00010_000101_00111; 
		615: oled_colour = 16'b00010_000101_00111; 
		616: oled_colour = 16'b00010_000101_00111; 
		617: oled_colour = 16'b00010_000101_00111; 
		618: oled_colour = 16'b00010_000101_00111; 
		619: oled_colour = 16'b00010_000101_00111; 
		620: oled_colour = 16'b00010_000101_00111; 
		621: oled_colour = 16'b00010_000101_00111; 
		622: oled_colour = 16'b00010_000101_00111; 
		623: oled_colour = 16'b00010_000101_00111; 
		624: oled_colour = 16'b00010_000101_00111; 
		625: oled_colour = 16'b00010_000101_00111; 
		626: oled_colour = 16'b00011_000101_00111; 
		627: oled_colour = 16'b00010_000101_00111; 
		628: oled_colour = 16'b00010_000101_00111; 
		629: oled_colour = 16'b00010_000101_00111; 
		630: oled_colour = 16'b00010_000101_00111; 
		631: oled_colour = 16'b00010_000101_00111; 
		632: oled_colour = 16'b00010_000101_00111; 
		633: oled_colour = 16'b00010_000101_00111; 
		634: oled_colour = 16'b00010_000101_00111; 
		635: oled_colour = 16'b00010_000101_00111; 
		636: oled_colour = 16'b00010_000101_00111; 
		637: oled_colour = 16'b00010_000101_01001; 
		638: oled_colour = 16'b00010_000111_01011; 
		639: oled_colour = 16'b00011_001100_01101; 
		640: oled_colour = 16'b00101_010001_01110; 
		641: oled_colour = 16'b00111_010101_01111; 
		642: oled_colour = 16'b01001_010111_10001; 
		643: oled_colour = 16'b01010_011010_10010; 
		644: oled_colour = 16'b01010_011010_10010; 
		645: oled_colour = 16'b01010_011010_10010; 
		646: oled_colour = 16'b01010_011001_10001; 
		647: oled_colour = 16'b01010_011001_10010; 
		648: oled_colour = 16'b01011_011010_10010; 
		649: oled_colour = 16'b01011_011010_10010; 
		650: oled_colour = 16'b01011_011011_10010; 
		651: oled_colour = 16'b01011_011011_10010; 
		652: oled_colour = 16'b01010_011001_10010; 
		653: oled_colour = 16'b01010_011001_10001; 
		654: oled_colour = 16'b01010_011010_10010; 
		655: oled_colour = 16'b01011_011010_10010; 
		656: oled_colour = 16'b01011_011011_10010; 
		657: oled_colour = 16'b01011_011011_10011; 
		658: oled_colour = 16'b01010_011010_10010; 
		659: oled_colour = 16'b01010_011001_10001; 
		660: oled_colour = 16'b01010_011001_10010; 
		661: oled_colour = 16'b01010_011000_10001; 
		662: oled_colour = 16'b01000_010100_01110; 
		663: oled_colour = 16'b00110_001111_01011; 
		664: oled_colour = 16'b01001_010100_01011; 
		665: oled_colour = 16'b01110_011111_01110; 
		666: oled_colour = 16'b01111_011111_01110; 
		667: oled_colour = 16'b10101_101010_10001; 
		668: oled_colour = 16'b10000_100010_01111; 
		669: oled_colour = 16'b10001_100011_10000; 
		670: oled_colour = 16'b10011_100111_10001; 
		671: oled_colour = 16'b01101_011101_01111; 
		672: oled_colour = 16'b01000_010110_10000; 
		673: oled_colour = 16'b01001_010111_10001; 
		674: oled_colour = 16'b01000_010101_10000; 
		675: oled_colour = 16'b00110_010011_01111; 
		676: oled_colour = 16'b00101_010001_01110; 
		677: oled_colour = 16'b00101_010000_01110; 
		678: oled_colour = 16'b00100_001111_01110; 
		679: oled_colour = 16'b00100_001101_01101; 
		680: oled_colour = 16'b00011_001011_01100; 
		681: oled_colour = 16'b00010_001001_01100; 
		682: oled_colour = 16'b00010_001001_01011; 
		683: oled_colour = 16'b00010_001001_01011; 
		684: oled_colour = 16'b00011_001010_01100; 
		685: oled_colour = 16'b00100_001011_01100; 
		686: oled_colour = 16'b00100_001110_01101; 
		687: oled_colour = 16'b00101_010000_01110; 
		688: oled_colour = 16'b00101_010000_01110; 
		689: oled_colour = 16'b00101_010000_01110; 
		690: oled_colour = 16'b00101_010000_01101; 
		691: oled_colour = 16'b00100_001111_01101; 
		692: oled_colour = 16'b00101_010000_01110; 
		693: oled_colour = 16'b00110_010001_01110; 
		694: oled_colour = 16'b00101_010010_01110; 
		695: oled_colour = 16'b00110_010010_01110; 
		696: oled_colour = 16'b00100_001111_01101; 
		697: oled_colour = 16'b00010_001001_01100; 
		698: oled_colour = 16'b00001_000100_01100; 
		699: oled_colour = 16'b01001_010101_01101; 
		700: oled_colour = 16'b11010_110000_01010; 
		701: oled_colour = 16'b11111_111011_00100; 
		702: oled_colour = 16'b11111_110110_01000; 
		703: oled_colour = 16'b01011_011001_01111; 
		704: oled_colour = 16'b00001_000111_01100; 
		705: oled_colour = 16'b00010_000100_01001; 
		706: oled_colour = 16'b00010_000101_01001; 
		707: oled_colour = 16'b00010_000101_01010; 
		708: oled_colour = 16'b00010_000100_01000; 
		709: oled_colour = 16'b00010_000101_00111; 
		710: oled_colour = 16'b00011_000101_00111; 
		711: oled_colour = 16'b00010_000101_00111; 
		712: oled_colour = 16'b00010_000101_00111; 
		713: oled_colour = 16'b00010_000101_00111; 
		714: oled_colour = 16'b00010_000101_00111; 
		715: oled_colour = 16'b00010_000101_00111; 
		716: oled_colour = 16'b00010_000101_00111; 
		717: oled_colour = 16'b00010_000101_00111; 
		718: oled_colour = 16'b00010_000101_00111; 
		719: oled_colour = 16'b00011_000101_01000; 
		720: oled_colour = 16'b00011_000101_01000; 
		721: oled_colour = 16'b00010_000101_01000; 
		722: oled_colour = 16'b00011_000101_01001; 
		723: oled_colour = 16'b00011_000101_01001; 
		724: oled_colour = 16'b00011_000101_01001; 
		725: oled_colour = 16'b00010_000101_01000; 
		726: oled_colour = 16'b00010_000101_01000; 
		727: oled_colour = 16'b00011_000101_01000; 
		728: oled_colour = 16'b00010_000101_00111; 
		729: oled_colour = 16'b00010_000101_00111; 
		730: oled_colour = 16'b00010_000101_00111; 
		731: oled_colour = 16'b00010_000101_00111; 
		732: oled_colour = 16'b00010_000101_00111; 
		733: oled_colour = 16'b00010_000101_01000; 
		734: oled_colour = 16'b00010_000110_01010; 
		735: oled_colour = 16'b00011_001000_01011; 
		736: oled_colour = 16'b00011_001100_01101; 
		737: oled_colour = 16'b00100_001110_01101; 
		738: oled_colour = 16'b00101_010000_01110; 
		739: oled_colour = 16'b00110_010001_01111; 
		740: oled_colour = 16'b00101_010000_01110; 
		741: oled_colour = 16'b00100_001110_01101; 
		742: oled_colour = 16'b00101_001111_01110; 
		743: oled_colour = 16'b00101_010001_01111; 
		744: oled_colour = 16'b00101_010000_01110; 
		745: oled_colour = 16'b00110_010010_01111; 
		746: oled_colour = 16'b00110_010010_01111; 
		747: oled_colour = 16'b00110_010001_01111; 
		748: oled_colour = 16'b00110_010010_01111; 
		749: oled_colour = 16'b00101_010001_01110; 
		750: oled_colour = 16'b00101_010000_01110; 
		751: oled_colour = 16'b00110_010010_01111; 
		752: oled_colour = 16'b00110_010010_01111; 
		753: oled_colour = 16'b00110_010001_01111; 
		754: oled_colour = 16'b00110_010010_01111; 
		755: oled_colour = 16'b00110_010010_01111; 
		756: oled_colour = 16'b00111_010100_10000; 
		757: oled_colour = 16'b01000_010101_10000; 
		758: oled_colour = 16'b01001_010111_10001; 
		759: oled_colour = 16'b01010_011001_10001; 
		760: oled_colour = 16'b00110_001111_01100; 
		761: oled_colour = 16'b00011_001010_01000; 
		762: oled_colour = 16'b00101_001101_01001; 
		763: oled_colour = 16'b00111_010000_01001; 
		764: oled_colour = 16'b01000_010010_01010; 
		765: oled_colour = 16'b01000_010001_01010; 
		766: oled_colour = 16'b01010_010110_01011; 
		767: oled_colour = 16'b01011_010111_01011; 
		768: oled_colour = 16'b01010_011001_10001; 
		769: oled_colour = 16'b01010_011001_10010; 
		770: oled_colour = 16'b01011_011001_10010; 
		771: oled_colour = 16'b01011_011010_10010; 
		772: oled_colour = 16'b01011_011010_10010; 
		773: oled_colour = 16'b01011_011010_10010; 
		774: oled_colour = 16'b01010_011010_10010; 
		775: oled_colour = 16'b01010_011001_10010; 
		776: oled_colour = 16'b01010_011001_10010; 
		777: oled_colour = 16'b01001_011000_10001; 
		778: oled_colour = 16'b01001_011000_10001; 
		779: oled_colour = 16'b01001_011000_10001; 
		780: oled_colour = 16'b01010_011001_10010; 
		781: oled_colour = 16'b01011_011010_10010; 
		782: oled_colour = 16'b01011_011011_10011; 
		783: oled_colour = 16'b01011_011010_10010; 
		784: oled_colour = 16'b01010_011001_10010; 
		785: oled_colour = 16'b01001_010111_10001; 
		786: oled_colour = 16'b00111_010101_10000; 
		787: oled_colour = 16'b00101_010001_01110; 
		788: oled_colour = 16'b00100_001101_01101; 
		789: oled_colour = 16'b00011_001010_01100; 
		790: oled_colour = 16'b00011_001001_01011; 
		791: oled_colour = 16'b00100_001011_01100; 
		792: oled_colour = 16'b00111_001111_01100; 
		793: oled_colour = 16'b01010_010011_01011; 
		794: oled_colour = 16'b01101_011100_01100; 
		795: oled_colour = 16'b11110_110110_00111; 
		796: oled_colour = 16'b11111_111010_00011; 
		797: oled_colour = 16'b11111_111000_00100; 
		798: oled_colour = 16'b11010_101111_01001; 
		799: oled_colour = 16'b01011_010111_01110; 
		800: oled_colour = 16'b00111_001111_01101; 
		801: oled_colour = 16'b00101_001100_01100; 
		802: oled_colour = 16'b00100_001100_01100; 
		803: oled_colour = 16'b00101_001111_01110; 
		804: oled_colour = 16'b00100_001101_01101; 
		805: oled_colour = 16'b00011_001011_01100; 
		806: oled_colour = 16'b00010_000111_01011; 
		807: oled_colour = 16'b00010_000101_01001; 
		808: oled_colour = 16'b00011_000101_01000; 
		809: oled_colour = 16'b00010_000101_00111; 
		810: oled_colour = 16'b00010_000101_00111; 
		811: oled_colour = 16'b00011_000101_00111; 
		812: oled_colour = 16'b00011_000101_00111; 
		813: oled_colour = 16'b00011_000101_00111; 
		814: oled_colour = 16'b00011_000101_00111; 
		815: oled_colour = 16'b00011_000101_00111; 
		816: oled_colour = 16'b00011_000101_01000; 
		817: oled_colour = 16'b00011_000101_01000; 
		818: oled_colour = 16'b00011_000101_00111; 
		819: oled_colour = 16'b00011_000101_00111; 
		820: oled_colour = 16'b00011_000101_00111; 
		821: oled_colour = 16'b00011_000101_00111; 
		822: oled_colour = 16'b00010_000101_00111; 
		823: oled_colour = 16'b00010_000101_00111; 
		824: oled_colour = 16'b00010_000101_00111; 
		825: oled_colour = 16'b00010_000101_00111; 
		826: oled_colour = 16'b00010_000101_00111; 
		827: oled_colour = 16'b00010_000101_00111; 
		828: oled_colour = 16'b00010_000101_00111; 
		829: oled_colour = 16'b00011_000101_01000; 
		830: oled_colour = 16'b00010_000101_01000; 
		831: oled_colour = 16'b00010_000101_01000; 
		832: oled_colour = 16'b00010_000101_01001; 
		833: oled_colour = 16'b00010_000110_01001; 
		834: oled_colour = 16'b00010_000101_01001; 
		835: oled_colour = 16'b00010_000101_01000; 
		836: oled_colour = 16'b00010_000100_01000; 
		837: oled_colour = 16'b00010_000100_01001; 
		838: oled_colour = 16'b00010_000100_01001; 
		839: oled_colour = 16'b00010_000100_01001; 
		840: oled_colour = 16'b00001_000100_01001; 
		841: oled_colour = 16'b00001_000100_01001; 
		842: oled_colour = 16'b00010_000100_01001; 
		843: oled_colour = 16'b00010_000100_01001; 
		844: oled_colour = 16'b00001_000101_01010; 
		845: oled_colour = 16'b00001_000101_01001; 
		846: oled_colour = 16'b00001_000100_01001; 
		847: oled_colour = 16'b00010_000100_01001; 
		848: oled_colour = 16'b00010_000100_01001; 
		849: oled_colour = 16'b00001_000100_01001; 
		850: oled_colour = 16'b00001_000100_01010; 
		851: oled_colour = 16'b00010_000101_01010; 
		852: oled_colour = 16'b00010_000110_01010; 
		853: oled_colour = 16'b00011_001000_01011; 
		854: oled_colour = 16'b00010_001000_01011; 
		855: oled_colour = 16'b00011_001100_01101; 
		856: oled_colour = 16'b00101_001111_01011; 
		857: oled_colour = 16'b00100_001011_00111; 
		858: oled_colour = 16'b00110_001111_01010; 
		859: oled_colour = 16'b00110_001111_01001; 
		860: oled_colour = 16'b00110_001110_01001; 
		861: oled_colour = 16'b00110_001110_01001; 
		862: oled_colour = 16'b00101_001101_01001; 
		863: oled_colour = 16'b00110_001101_01001; 
		864: oled_colour = 16'b01100_011010_01110; 
		865: oled_colour = 16'b01000_010110_10001; 
		866: oled_colour = 16'b01001_011000_10001; 
		867: oled_colour = 16'b01001_011000_10001; 
		868: oled_colour = 16'b01001_011000_10001; 
		869: oled_colour = 16'b01001_011000_10001; 
		870: oled_colour = 16'b01010_011001_10010; 
		871: oled_colour = 16'b01010_011001_10010; 
		872: oled_colour = 16'b01010_011001_10010; 
		873: oled_colour = 16'b01011_011010_10010; 
		874: oled_colour = 16'b01011_011010_10010; 
		875: oled_colour = 16'b01010_011001_10010; 
		876: oled_colour = 16'b01010_011000_10010; 
		877: oled_colour = 16'b01001_010110_10001; 
		878: oled_colour = 16'b01001_010101_10001; 
		879: oled_colour = 16'b01001_010101_10001; 
		880: oled_colour = 16'b01000_010110_10001; 
		881: oled_colour = 16'b01001_011000_10001; 
		882: oled_colour = 16'b01001_011001_10001; 
		883: oled_colour = 16'b01010_011001_10010; 
		884: oled_colour = 16'b01010_011001_10010; 
		885: oled_colour = 16'b01010_011001_10010; 
		886: oled_colour = 16'b01010_011001_10010; 
		887: oled_colour = 16'b01100_011011_10011; 
		888: oled_colour = 16'b10000_100010_10011; 
		889: oled_colour = 16'b11001_101101_10001; 
		890: oled_colour = 16'b11101_110100_01100; 
		891: oled_colour = 16'b11100_110010_01010; 
		892: oled_colour = 16'b11011_110010_01011; 
		893: oled_colour = 16'b11011_110001_01011; 
		894: oled_colour = 16'b10101_101000_01111; 
		895: oled_colour = 16'b01111_100000_10010; 
		896: oled_colour = 16'b01010_011001_10001; 
		897: oled_colour = 16'b00111_010100_10000; 
		898: oled_colour = 16'b00110_010001_01111; 
		899: oled_colour = 16'b00101_001111_01110; 
		900: oled_colour = 16'b00101_001111_01110; 
		901: oled_colour = 16'b00011_001011_01100; 
		902: oled_colour = 16'b00010_000111_01011; 
		903: oled_colour = 16'b00010_000101_01010; 
		904: oled_colour = 16'b00010_000101_01001; 
		905: oled_colour = 16'b00010_000100_01001; 
		906: oled_colour = 16'b00010_000101_01001; 
		907: oled_colour = 16'b00010_000101_01001; 
		908: oled_colour = 16'b00010_000101_01001; 
		909: oled_colour = 16'b00010_000100_01001; 
		910: oled_colour = 16'b00010_000100_01001; 
		911: oled_colour = 16'b00010_000100_01001; 
		912: oled_colour = 16'b00010_000100_01000; 
		913: oled_colour = 16'b00010_000100_01000; 
		914: oled_colour = 16'b00010_000100_01000; 
		915: oled_colour = 16'b00010_000100_01000; 
		916: oled_colour = 16'b00010_000100_01000; 
		917: oled_colour = 16'b00010_000100_01000; 
		918: oled_colour = 16'b00010_000100_01000; 
		919: oled_colour = 16'b00010_000101_01000; 
		920: oled_colour = 16'b00011_000101_01001; 
		921: oled_colour = 16'b00010_000101_01001; 
		922: oled_colour = 16'b00011_000101_01000; 
		923: oled_colour = 16'b00011_000101_01000; 
		924: oled_colour = 16'b00011_000101_01000; 
		925: oled_colour = 16'b00011_000101_01000; 
		926: oled_colour = 16'b00011_000101_01000; 
		927: oled_colour = 16'b00010_000101_01000; 
		928: oled_colour = 16'b00011_000101_01000; 
		929: oled_colour = 16'b00010_000101_01000; 
		930: oled_colour = 16'b00010_000101_01001; 
		931: oled_colour = 16'b00010_000110_01010; 
		932: oled_colour = 16'b00011_001000_01011; 
		933: oled_colour = 16'b00100_001101_01101; 
		934: oled_colour = 16'b00110_010000_01110; 
		935: oled_colour = 16'b00110_010001_01110; 
		936: oled_colour = 16'b00110_010001_01110; 
		937: oled_colour = 16'b00110_010000_01110; 
		938: oled_colour = 16'b00110_001111_01110; 
		939: oled_colour = 16'b00110_001111_01110; 
		940: oled_colour = 16'b00110_010001_01111; 
		941: oled_colour = 16'b00110_010001_01111; 
		942: oled_colour = 16'b00110_010000_01110; 
		943: oled_colour = 16'b00110_010000_01110; 
		944: oled_colour = 16'b00110_001111_01110; 
		945: oled_colour = 16'b00101_001111_01110; 
		946: oled_colour = 16'b00110_010001_01110; 
		947: oled_colour = 16'b00111_010011_01111; 
		948: oled_colour = 16'b00111_010011_01111; 
		949: oled_colour = 16'b00110_010010_01111; 
		950: oled_colour = 16'b00110_010001_01111; 
		951: oled_colour = 16'b00110_010001_01111; 
		952: oled_colour = 16'b00101_001111_01011; 
		953: oled_colour = 16'b00011_001011_00111; 
		954: oled_colour = 16'b00110_001110_01001; 
		955: oled_colour = 16'b01101_011011_01101; 
		956: oled_colour = 16'b00101_001111_01001; 
		957: oled_colour = 16'b00111_001111_01001; 
		958: oled_colour = 16'b01011_011000_01011; 
		959: oled_colour = 16'b00111_010000_01001; 
		960: oled_colour = 16'b01011_010110_01011; 
		961: oled_colour = 16'b00011_001010_01100; 
		962: oled_colour = 16'b00100_001101_01101; 
		963: oled_colour = 16'b00011_001101_01101; 
		964: oled_colour = 16'b00100_001101_01101; 
		965: oled_colour = 16'b00100_001101_01101; 
		966: oled_colour = 16'b00100_001110_01101; 
		967: oled_colour = 16'b00100_001110_01101; 
		968: oled_colour = 16'b00100_010000_01110; 
		969: oled_colour = 16'b00101_010001_01110; 
		970: oled_colour = 16'b00101_010010_01111; 
		971: oled_colour = 16'b00101_010000_01110; 
		972: oled_colour = 16'b00100_001110_01101; 
		973: oled_colour = 16'b00011_001100_01101; 
		974: oled_colour = 16'b00010_001010_01101; 
		975: oled_colour = 16'b00010_001000_01100; 
		976: oled_colour = 16'b00010_001000_01100; 
		977: oled_colour = 16'b00011_001011_01100; 
		978: oled_colour = 16'b00100_001101_01101; 
		979: oled_colour = 16'b00100_001110_01101; 
		980: oled_colour = 16'b00101_010000_01110; 
		981: oled_colour = 16'b00110_010011_01111; 
		982: oled_colour = 16'b00111_010100_10000; 
		983: oled_colour = 16'b01010_010111_10000; 
		984: oled_colour = 16'b01110_011011_01110; 
		985: oled_colour = 16'b10010_100011_01101; 
		986: oled_colour = 16'b11111_110101_01000; 
		987: oled_colour = 16'b11111_111000_00101; 
		988: oled_colour = 16'b11111_111000_00100; 
		989: oled_colour = 16'b11110_110100_01001; 
		990: oled_colour = 16'b01111_011110_01111; 
		991: oled_colour = 16'b00101_001111_01110; 
		992: oled_colour = 16'b00011_001101_01101; 
		993: oled_colour = 16'b00010_001011_01100; 
		994: oled_colour = 16'b00010_001001_01100; 
		995: oled_colour = 16'b00011_000111_01011; 
		996: oled_colour = 16'b00011_001011_01100; 
		997: oled_colour = 16'b00011_001010_01100; 
		998: oled_colour = 16'b00100_001001_01100; 
		999: oled_colour = 16'b00100_001010_01100; 
		1000: oled_colour = 16'b00011_001010_01100; 
		1001: oled_colour = 16'b00011_001010_01100; 
		1002: oled_colour = 16'b00011_001011_01101; 
		1003: oled_colour = 16'b00100_001101_01101; 
		1004: oled_colour = 16'b00100_001101_01101; 
		1005: oled_colour = 16'b00100_001101_01101; 
		1006: oled_colour = 16'b00100_001101_01101; 
		1007: oled_colour = 16'b00101_001110_01110; 
		1008: oled_colour = 16'b00101_001111_01110; 
		1009: oled_colour = 16'b00101_001110_01110; 
		1010: oled_colour = 16'b00101_001110_01110; 
		1011: oled_colour = 16'b00110_010000_01110; 
		1012: oled_colour = 16'b00110_001111_01110; 
		1013: oled_colour = 16'b00101_001110_01110; 
		1014: oled_colour = 16'b00100_001101_01101; 
		1015: oled_colour = 16'b00011_001010_01100; 
		1016: oled_colour = 16'b00010_000111_01011; 
		1017: oled_colour = 16'b00010_000110_01011; 
		1018: oled_colour = 16'b00011_000110_01001; 
		1019: oled_colour = 16'b00011_000110_01001; 
		1020: oled_colour = 16'b00011_000110_01001; 
		1021: oled_colour = 16'b00011_000101_01001; 
		1022: oled_colour = 16'b00011_000101_01001; 
		1023: oled_colour = 16'b00011_000101_01001; 
		1024: oled_colour = 16'b00011_000101_01001; 
		1025: oled_colour = 16'b00011_000101_01001; 
		1026: oled_colour = 16'b00010_000110_01010; 
		1027: oled_colour = 16'b00010_000111_01100; 
		1028: oled_colour = 16'b00010_000111_01100; 
		1029: oled_colour = 16'b00011_001011_01101; 
		1030: oled_colour = 16'b00101_001101_01110; 
		1031: oled_colour = 16'b00101_001111_01110; 
		1032: oled_colour = 16'b00101_001110_01101; 
		1033: oled_colour = 16'b00100_001101_01101; 
		1034: oled_colour = 16'b00101_001110_01110; 
		1035: oled_colour = 16'b00100_001110_01110; 
		1036: oled_colour = 16'b00101_001110_01110; 
		1037: oled_colour = 16'b00101_001111_01110; 
		1038: oled_colour = 16'b00101_001110_01110; 
		1039: oled_colour = 16'b00100_001101_01101; 
		1040: oled_colour = 16'b00100_001110_01110; 
		1041: oled_colour = 16'b00100_001110_01101; 
		1042: oled_colour = 16'b00101_001110_01101; 
		1043: oled_colour = 16'b00101_001111_01110; 
		1044: oled_colour = 16'b00101_001111_01101; 
		1045: oled_colour = 16'b01010_011000_10000; 
		1046: oled_colour = 16'b01111_100000_10010; 
		1047: oled_colour = 16'b01111_100001_10010; 
		1048: oled_colour = 16'b01010_010110_01100; 
		1049: oled_colour = 16'b01001_010101_01011; 
		1050: oled_colour = 16'b01000_010011_01010; 
		1051: oled_colour = 16'b10001_100010_01111; 
		1052: oled_colour = 16'b00101_001111_01000; 
		1053: oled_colour = 16'b00101_001110_01000; 
		1054: oled_colour = 16'b10010_100100_01111; 
		1055: oled_colour = 16'b00101_001111_01000; 
		1056: oled_colour = 16'b01110_011010_01010; 
		1057: oled_colour = 16'b00011_000101_01000; 
		1058: oled_colour = 16'b00010_000101_01001; 
		1059: oled_colour = 16'b00010_000101_01001; 
		1060: oled_colour = 16'b00010_000101_01001; 
		1061: oled_colour = 16'b00010_000101_01001; 
		1062: oled_colour = 16'b00010_000101_01001; 
		1063: oled_colour = 16'b00010_000101_01001; 
		1064: oled_colour = 16'b00010_000110_01010; 
		1065: oled_colour = 16'b00010_000110_01010; 
		1066: oled_colour = 16'b00010_000110_01010; 
		1067: oled_colour = 16'b00010_000110_01010; 
		1068: oled_colour = 16'b00010_000110_01010; 
		1069: oled_colour = 16'b00011_000110_01010; 
		1070: oled_colour = 16'b00011_000110_01010; 
		1071: oled_colour = 16'b00011_000110_01010; 
		1072: oled_colour = 16'b00011_000101_01001; 
		1073: oled_colour = 16'b00011_000101_01001; 
		1074: oled_colour = 16'b00010_000101_01010; 
		1075: oled_colour = 16'b00010_000110_01010; 
		1076: oled_colour = 16'b00010_000101_01010; 
		1077: oled_colour = 16'b00010_000101_01001; 
		1078: oled_colour = 16'b00010_000101_01001; 
		1079: oled_colour = 16'b00010_000100_01000; 
		1080: oled_colour = 16'b00001_000001_01001; 
		1081: oled_colour = 16'b01001_010100_01111; 
		1082: oled_colour = 16'b11111_111011_00100; 
		1083: oled_colour = 16'b11111_111100_00001; 
		1084: oled_colour = 16'b11111_111001_00011; 
		1085: oled_colour = 16'b11100_110001_01010; 
		1086: oled_colour = 16'b01001_010110_01111; 
		1087: oled_colour = 16'b00001_001001_01100; 
		1088: oled_colour = 16'b00100_001101_01101; 
		1089: oled_colour = 16'b00111_010010_01111; 
		1090: oled_colour = 16'b01000_010101_10000; 
		1091: oled_colour = 16'b01000_010101_10000; 
		1092: oled_colour = 16'b01000_010101_10000; 
		1093: oled_colour = 16'b01000_010110_10001; 
		1094: oled_colour = 16'b01010_011001_10010; 
		1095: oled_colour = 16'b01011_011011_10010; 
		1096: oled_colour = 16'b01100_011100_10010; 
		1097: oled_colour = 16'b01011_011011_10010; 
		1098: oled_colour = 16'b01100_011100_10010; 
		1099: oled_colour = 16'b01100_011100_10010; 
		1100: oled_colour = 16'b01100_011100_10010; 
		1101: oled_colour = 16'b01100_011100_10010; 
		1102: oled_colour = 16'b01011_011011_10010; 
		1103: oled_colour = 16'b01011_011100_10010; 
		1104: oled_colour = 16'b01011_011011_10010; 
		1105: oled_colour = 16'b01011_011010_10001; 
		1106: oled_colour = 16'b01011_011010_10001; 
		1107: oled_colour = 16'b01010_011000_10001; 
		1108: oled_colour = 16'b01001_010110_10001; 
		1109: oled_colour = 16'b01000_010100_10000; 
		1110: oled_colour = 16'b00111_010010_01111; 
		1111: oled_colour = 16'b00100_001110_01101; 
		1112: oled_colour = 16'b00011_000111_01011; 
		1113: oled_colour = 16'b00011_000101_01001; 
		1114: oled_colour = 16'b00011_000110_01001; 
		1115: oled_colour = 16'b00011_000101_01001; 
		1116: oled_colour = 16'b00011_000101_01001; 
		1117: oled_colour = 16'b00011_000101_01001; 
		1118: oled_colour = 16'b00011_000101_01001; 
		1119: oled_colour = 16'b00011_000101_01001; 
		1120: oled_colour = 16'b00011_000101_01001; 
		1121: oled_colour = 16'b00011_000101_01001; 
		1122: oled_colour = 16'b00011_000110_01001; 
		1123: oled_colour = 16'b00011_000101_01001; 
		1124: oled_colour = 16'b00011_000101_01001; 
		1125: oled_colour = 16'b00010_000100_01001; 
		1126: oled_colour = 16'b00010_000100_01001; 
		1127: oled_colour = 16'b00010_000100_01001; 
		1128: oled_colour = 16'b00010_000100_01001; 
		1129: oled_colour = 16'b00010_000100_01001; 
		1130: oled_colour = 16'b00010_000101_01001; 
		1131: oled_colour = 16'b00010_000100_01001; 
		1132: oled_colour = 16'b00010_000100_01001; 
		1133: oled_colour = 16'b00010_000100_01001; 
		1134: oled_colour = 16'b00010_000100_01001; 
		1135: oled_colour = 16'b00010_000100_01001; 
		1136: oled_colour = 16'b00010_000100_01001; 
		1137: oled_colour = 16'b00010_000100_01001; 
		1138: oled_colour = 16'b00010_000100_01001; 
		1139: oled_colour = 16'b00001_000011_01000; 
		1140: oled_colour = 16'b00110_001101_01100; 
		1141: oled_colour = 16'b01100_011001_01110; 
		1142: oled_colour = 16'b01100_011010_01101; 
		1143: oled_colour = 16'b01001_010100_01011; 
		1144: oled_colour = 16'b01001_010011_01011; 
		1145: oled_colour = 16'b01000_010001_01010; 
		1146: oled_colour = 16'b00110_001101_01001; 
		1147: oled_colour = 16'b10000_100001_01111; 
		1148: oled_colour = 16'b01001_010101_01010; 
		1149: oled_colour = 16'b00101_001101_01000; 
		1150: oled_colour = 16'b10000_100000_01110; 
		1151: oled_colour = 16'b01010_010110_01011; 
		1152: oled_colour = 16'b01111_011101_01010; 
		1153: oled_colour = 16'b01000_001111_01001; 
		1154: oled_colour = 16'b00010_000100_01010; 
		1155: oled_colour = 16'b00011_000110_01010; 
		1156: oled_colour = 16'b00011_000110_01010; 
		1157: oled_colour = 16'b00011_000110_01010; 
		1158: oled_colour = 16'b00011_000110_01010; 
		1159: oled_colour = 16'b00011_000110_01010; 
		1160: oled_colour = 16'b00011_000110_01010; 
		1161: oled_colour = 16'b00011_000110_01010; 
		1162: oled_colour = 16'b00011_000101_01001; 
		1163: oled_colour = 16'b00011_000101_01001; 
		1164: oled_colour = 16'b00011_000101_01001; 
		1165: oled_colour = 16'b00011_000101_01001; 
		1166: oled_colour = 16'b00011_000101_01001; 
		1167: oled_colour = 16'b00011_000101_01001; 
		1168: oled_colour = 16'b00011_000101_01001; 
		1169: oled_colour = 16'b00010_000101_01001; 
		1170: oled_colour = 16'b00010_000100_01001; 
		1171: oled_colour = 16'b00010_000100_01001; 
		1172: oled_colour = 16'b00010_000100_01001; 
		1173: oled_colour = 16'b00010_000101_01001; 
		1174: oled_colour = 16'b00011_001000_01010; 
		1175: oled_colour = 16'b00110_001100_01100; 
		1176: oled_colour = 16'b01001_010011_01101; 
		1177: oled_colour = 16'b10101_101000_01011; 
		1178: oled_colour = 16'b11111_111011_00011; 
		1179: oled_colour = 16'b11111_111010_00001; 
		1180: oled_colour = 16'b11111_111010_00010; 
		1181: oled_colour = 16'b11111_110101_00111; 
		1182: oled_colour = 16'b10010_100100_01110; 
		1183: oled_colour = 16'b01001_010101_01110; 
		1184: oled_colour = 16'b00111_010000_01110; 
		1185: oled_colour = 16'b00101_001110_01101; 
		1186: oled_colour = 16'b00100_001100_01101; 
		1187: oled_colour = 16'b00101_001111_01110; 
		1188: oled_colour = 16'b00110_010001_01111; 
		1189: oled_colour = 16'b00111_010100_01111; 
		1190: oled_colour = 16'b01011_011010_10001; 
		1191: oled_colour = 16'b01101_011101_10010; 
		1192: oled_colour = 16'b01101_011101_10010; 
		1193: oled_colour = 16'b01101_011110_10010; 
		1194: oled_colour = 16'b01101_011110_10010; 
		1195: oled_colour = 16'b01101_011110_10010; 
		1196: oled_colour = 16'b01101_011101_10010; 
		1197: oled_colour = 16'b01101_011100_10010; 
		1198: oled_colour = 16'b01010_011000_10001; 
		1199: oled_colour = 16'b00110_010001_01110; 
		1200: oled_colour = 16'b00100_001110_01101; 
		1201: oled_colour = 16'b00011_001011_01100; 
		1202: oled_colour = 16'b00011_001001_01100; 
		1203: oled_colour = 16'b00010_001000_01011; 
		1204: oled_colour = 16'b00010_000111_01011; 
		1205: oled_colour = 16'b00010_000110_01011; 
		1206: oled_colour = 16'b00001_000101_01011; 
		1207: oled_colour = 16'b00010_000101_01010; 
		1208: oled_colour = 16'b00010_000101_01010; 
		1209: oled_colour = 16'b00010_000101_01010; 
		1210: oled_colour = 16'b00001_000101_01010; 
		1211: oled_colour = 16'b00010_000101_01010; 
		1212: oled_colour = 16'b00010_000101_01010; 
		1213: oled_colour = 16'b00011_000110_01010; 
		1214: oled_colour = 16'b00011_000101_01001; 
		1215: oled_colour = 16'b00011_000110_01001; 
		1216: oled_colour = 16'b00011_000101_01001; 
		1217: oled_colour = 16'b00011_000101_01001; 
		1218: oled_colour = 16'b00011_000101_01001; 
		1219: oled_colour = 16'b00011_000101_01001; 
		1220: oled_colour = 16'b00011_000101_01001; 
		1221: oled_colour = 16'b00011_000110_01001; 
		1222: oled_colour = 16'b00011_000110_01001; 
		1223: oled_colour = 16'b00011_000110_01001; 
		1224: oled_colour = 16'b00011_000110_01001; 
		1225: oled_colour = 16'b00011_000110_01001; 
		1226: oled_colour = 16'b00011_000110_01001; 
		1227: oled_colour = 16'b00011_000110_01001; 
		1228: oled_colour = 16'b00011_000110_01001; 
		1229: oled_colour = 16'b00011_000110_01001; 
		1230: oled_colour = 16'b00011_000110_01001; 
		1231: oled_colour = 16'b00011_000110_01001; 
		1232: oled_colour = 16'b00011_000110_01001; 
		1233: oled_colour = 16'b00011_000110_01001; 
		1234: oled_colour = 16'b00011_000110_01001; 
		1235: oled_colour = 16'b00011_000101_01001; 
		1236: oled_colour = 16'b00101_001010_01010; 
		1237: oled_colour = 16'b00101_001100_00111; 
		1238: oled_colour = 16'b00101_001110_01000; 
		1239: oled_colour = 16'b00111_010000_01001; 
		1240: oled_colour = 16'b01000_010011_01010; 
		1241: oled_colour = 16'b01011_011000_01011; 
		1242: oled_colour = 16'b00111_010001_01001; 
		1243: oled_colour = 16'b10000_100001_01110; 
		1244: oled_colour = 16'b01100_011001_01100; 
		1245: oled_colour = 16'b00011_001010_00111; 
		1246: oled_colour = 16'b10001_100010_01111; 
		1247: oled_colour = 16'b01100_011010_01100; 
		1248: oled_colour = 16'b01101_011010_01010; 
		1249: oled_colour = 16'b01110_011011_01010; 
		1250: oled_colour = 16'b00010_000101_01010; 
		1251: oled_colour = 16'b00011_000110_01010; 
		1252: oled_colour = 16'b00010_000101_01010; 
		1253: oled_colour = 16'b00010_000110_01010; 
		1254: oled_colour = 16'b00011_000110_01010; 
		1255: oled_colour = 16'b00010_000110_01001; 
		1256: oled_colour = 16'b00011_000110_01001; 
		1257: oled_colour = 16'b00011_000110_01001; 
		1258: oled_colour = 16'b00011_000110_01001; 
		1259: oled_colour = 16'b00011_000110_01001; 
		1260: oled_colour = 16'b00011_000101_01001; 
		1261: oled_colour = 16'b00011_000101_01001; 
		1262: oled_colour = 16'b00011_000101_01001; 
		1263: oled_colour = 16'b00011_000101_01010; 
		1264: oled_colour = 16'b00010_000110_01011; 
		1265: oled_colour = 16'b00011_001001_01100; 
		1266: oled_colour = 16'b00100_001101_01110; 
		1267: oled_colour = 16'b00101_010000_01110; 
		1268: oled_colour = 16'b00111_010011_01111; 
		1269: oled_colour = 16'b01001_010111_10001; 
		1270: oled_colour = 16'b01010_011001_10001; 
		1271: oled_colour = 16'b01101_011101_10010; 
		1272: oled_colour = 16'b10010_100100_10010; 
		1273: oled_colour = 16'b11000_101100_01111; 
		1274: oled_colour = 16'b11011_110000_01100; 
		1275: oled_colour = 16'b11100_110011_01010; 
		1276: oled_colour = 16'b11100_110011_01010; 
		1277: oled_colour = 16'b11010_110000_01100; 
		1278: oled_colour = 16'b10100_100110_10000; 
		1279: oled_colour = 16'b01110_011101_10010; 
		1280: oled_colour = 16'b01101_011101_10010; 
		1281: oled_colour = 16'b01100_011101_10010; 
		1282: oled_colour = 16'b01011_011011_10010; 
		1283: oled_colour = 16'b01100_011101_10010; 
		1284: oled_colour = 16'b01101_011110_10011; 
		1285: oled_colour = 16'b01101_011110_10010; 
		1286: oled_colour = 16'b01101_011110_10010; 
		1287: oled_colour = 16'b01100_011100_10010; 
		1288: oled_colour = 16'b01100_011011_10010; 
		1289: oled_colour = 16'b01011_011010_10001; 
		1290: oled_colour = 16'b01010_011000_10001; 
		1291: oled_colour = 16'b01010_011001_10001; 
		1292: oled_colour = 16'b01010_011001_10001; 
		1293: oled_colour = 16'b01010_011000_10000; 
		1294: oled_colour = 16'b01001_010111_10000; 
		1295: oled_colour = 16'b01010_011001_10001; 
		1296: oled_colour = 16'b01011_011010_10001; 
		1297: oled_colour = 16'b01011_011010_10001; 
		1298: oled_colour = 16'b01010_011001_10001; 
		1299: oled_colour = 16'b01010_011000_10001; 
		1300: oled_colour = 16'b01001_010111_10001; 
		1301: oled_colour = 16'b01001_010111_10001; 
		1302: oled_colour = 16'b01001_010111_10001; 
		1303: oled_colour = 16'b01000_010110_10000; 
		1304: oled_colour = 16'b01000_010100_10000; 
		1305: oled_colour = 16'b00111_010011_10000; 
		1306: oled_colour = 16'b00110_010011_01111; 
		1307: oled_colour = 16'b00110_010010_01111; 
		1308: oled_colour = 16'b00110_010001_01111; 
		1309: oled_colour = 16'b00100_001111_01110; 
		1310: oled_colour = 16'b00010_001001_01100; 
		1311: oled_colour = 16'b00010_000110_01011; 
		1312: oled_colour = 16'b00011_000101_01010; 
		1313: oled_colour = 16'b00011_000101_01001; 
		1314: oled_colour = 16'b00011_000101_01001; 
		1315: oled_colour = 16'b00011_000101_01001; 
		1316: oled_colour = 16'b00011_000101_01001; 
		1317: oled_colour = 16'b00011_000101_01001; 
		1318: oled_colour = 16'b00011_000101_01001; 
		1319: oled_colour = 16'b00011_000101_01001; 
		1320: oled_colour = 16'b00011_000101_01001; 
		1321: oled_colour = 16'b00011_000101_01001; 
		1322: oled_colour = 16'b00011_000101_01001; 
		1323: oled_colour = 16'b00011_000101_01001; 
		1324: oled_colour = 16'b00011_000101_01001; 
		1325: oled_colour = 16'b00011_000101_01001; 
		1326: oled_colour = 16'b00011_000101_01001; 
		1327: oled_colour = 16'b00011_000101_01001; 
		1328: oled_colour = 16'b00011_000101_01001; 
		1329: oled_colour = 16'b00011_000101_01001; 
		1330: oled_colour = 16'b00011_000101_01001; 
		1331: oled_colour = 16'b00011_000110_01001; 
		1332: oled_colour = 16'b00111_001110_01011; 
		1333: oled_colour = 16'b00111_010000_01000; 
		1334: oled_colour = 16'b01101_011101_01110; 
		1335: oled_colour = 16'b01100_011011_01101; 
		1336: oled_colour = 16'b01011_011000_01100; 
		1337: oled_colour = 16'b01001_010100_01011; 
		1338: oled_colour = 16'b00100_001100_01000; 
		1339: oled_colour = 16'b01101_011010_01101; 
		1340: oled_colour = 16'b01101_011010_01100; 
		1341: oled_colour = 16'b00100_001010_01000; 
		1342: oled_colour = 16'b01101_011011_01101; 
		1343: oled_colour = 16'b01101_011011_01100; 
		1344: oled_colour = 16'b01100_010111_01010; 
		1345: oled_colour = 16'b10000_011110_01010; 
		1346: oled_colour = 16'b01000_001110_01000; 
		1347: oled_colour = 16'b00001_000011_01000; 
		1348: oled_colour = 16'b00011_000110_01001; 
		1349: oled_colour = 16'b00011_000101_01001; 
		1350: oled_colour = 16'b00011_000101_01001; 
		1351: oled_colour = 16'b00011_000101_01001; 
		1352: oled_colour = 16'b00011_000101_01001; 
		1353: oled_colour = 16'b00011_000101_01001; 
		1354: oled_colour = 16'b00011_000101_01001; 
		1355: oled_colour = 16'b00011_000101_01001; 
		1356: oled_colour = 16'b00011_000101_01001; 
		1357: oled_colour = 16'b00011_000101_01001; 
		1358: oled_colour = 16'b00011_000110_01001; 
		1359: oled_colour = 16'b00011_000101_01001; 
		1360: oled_colour = 16'b00011_000111_01011; 
		1361: oled_colour = 16'b00100_001100_01101; 
		1362: oled_colour = 16'b00110_010001_01111; 
		1363: oled_colour = 16'b00111_010011_01111; 
		1364: oled_colour = 16'b00111_010010_01111; 
		1365: oled_colour = 16'b00111_010010_01111; 
		1366: oled_colour = 16'b00111_010100_01111; 
		1367: oled_colour = 16'b01010_011000_10000; 
		1368: oled_colour = 16'b01110_011110_10001; 
		1369: oled_colour = 16'b10110_101001_01111; 
		1370: oled_colour = 16'b11110_110101_01001; 
		1371: oled_colour = 16'b11110_110101_00111; 
		1372: oled_colour = 16'b11101_110101_01000; 
		1373: oled_colour = 16'b11100_110011_01001; 
		1374: oled_colour = 16'b11010_101111_01100; 
		1375: oled_colour = 16'b10100_100110_01111; 
		1376: oled_colour = 16'b01101_011100_10001; 
		1377: oled_colour = 16'b01010_010111_10001; 
		1378: oled_colour = 16'b01000_010101_10000; 
		1379: oled_colour = 16'b00110_010010_01111; 
		1380: oled_colour = 16'b00101_010001_01110; 
		1381: oled_colour = 16'b00101_001111_01101; 
		1382: oled_colour = 16'b00100_001101_01101; 
		1383: oled_colour = 16'b00011_001101_01101; 
		1384: oled_colour = 16'b00101_010000_01110; 
		1385: oled_colour = 16'b00110_010010_01110; 
		1386: oled_colour = 16'b01000_010110_10000; 
		1387: oled_colour = 16'b01001_011000_10001; 
		1388: oled_colour = 16'b01011_011010_10010; 
		1389: oled_colour = 16'b01011_011011_10010; 
		1390: oled_colour = 16'b01011_011011_10001; 
		1391: oled_colour = 16'b01100_011100_10010; 
		1392: oled_colour = 16'b01101_011101_10010; 
		1393: oled_colour = 16'b01101_011110_10011; 
		1394: oled_colour = 16'b01101_011101_10010; 
		1395: oled_colour = 16'b01100_011100_10010; 
		1396: oled_colour = 16'b01011_011011_10010; 
		1397: oled_colour = 16'b01001_010111_10001; 
		1398: oled_colour = 16'b00110_010011_01111; 
		1399: oled_colour = 16'b00110_010010_01110; 
		1400: oled_colour = 16'b00110_010000_01110; 
		1401: oled_colour = 16'b00101_001111_01110; 
		1402: oled_colour = 16'b00101_001111_01110; 
		1403: oled_colour = 16'b00100_001101_01101; 
		1404: oled_colour = 16'b00011_001010_01100; 
		1405: oled_colour = 16'b00011_001000_01011; 
		1406: oled_colour = 16'b00010_000111_01010; 
		1407: oled_colour = 16'b00010_000110_01010; 
		1408: oled_colour = 16'b00011_000101_01001; 
		1409: oled_colour = 16'b00011_000101_01001; 
		1410: oled_colour = 16'b00011_000101_01001; 
		1411: oled_colour = 16'b00011_000101_01001; 
		1412: oled_colour = 16'b00011_000101_01001; 
		1413: oled_colour = 16'b00011_000101_01001; 
		1414: oled_colour = 16'b00011_000101_01001; 
		1415: oled_colour = 16'b00011_000101_01001; 
		1416: oled_colour = 16'b00011_000101_01001; 
		1417: oled_colour = 16'b00011_000101_01001; 
		1418: oled_colour = 16'b00011_000101_01001; 
		1419: oled_colour = 16'b00011_000101_01001; 
		1420: oled_colour = 16'b00011_000101_01001; 
		1421: oled_colour = 16'b00011_000101_01001; 
		1422: oled_colour = 16'b00011_000101_01001; 
		1423: oled_colour = 16'b00011_000101_01001; 
		1424: oled_colour = 16'b00011_000101_01001; 
		1425: oled_colour = 16'b00011_000101_01001; 
		1426: oled_colour = 16'b00011_000101_01001; 
		1427: oled_colour = 16'b00011_000111_01010; 
		1428: oled_colour = 16'b01000_010000_01011; 
		1429: oled_colour = 16'b00101_001010_00110; 
		1430: oled_colour = 16'b00100_001010_01000; 
		1431: oled_colour = 16'b00100_001001_00111; 
		1432: oled_colour = 16'b00101_001110_01000; 
		1433: oled_colour = 16'b00111_010010_01001; 
		1434: oled_colour = 16'b00110_010000_01001; 
		1435: oled_colour = 16'b01110_011100_01101; 
		1436: oled_colour = 16'b10000_100010_01110; 
		1437: oled_colour = 16'b00011_001010_00111; 
		1438: oled_colour = 16'b01100_011001_01101; 
		1439: oled_colour = 16'b10001_100011_01111; 
		1440: oled_colour = 16'b01011_010110_01010; 
		1441: oled_colour = 16'b01110_011011_01010; 
		1442: oled_colour = 16'b01111_011011_01010; 
		1443: oled_colour = 16'b00010_000100_01001; 
		1444: oled_colour = 16'b00011_000110_01010; 
		1445: oled_colour = 16'b00010_000110_01011; 
		1446: oled_colour = 16'b00010_000111_01100; 
		1447: oled_colour = 16'b00010_001001_01100; 
		1448: oled_colour = 16'b00010_001010_01100; 
		1449: oled_colour = 16'b00010_001000_01100; 
		1450: oled_colour = 16'b00010_000110_01011; 
		1451: oled_colour = 16'b00010_000110_01010; 
		1452: oled_colour = 16'b00011_000110_01010; 
		1453: oled_colour = 16'b00011_000101_01010; 
		1454: oled_colour = 16'b00011_000101_01010; 
		1455: oled_colour = 16'b00010_000101_01010; 
		1456: oled_colour = 16'b00010_000101_01010; 
		1457: oled_colour = 16'b00010_000100_01001; 
		1458: oled_colour = 16'b00010_000101_01010; 
		1459: oled_colour = 16'b00010_000101_01010; 
		1460: oled_colour = 16'b00010_000101_01011; 
		1461: oled_colour = 16'b00010_000101_01011; 
		1462: oled_colour = 16'b00010_000101_01011; 
		1463: oled_colour = 16'b00010_000110_01011; 
		1464: oled_colour = 16'b00100_001001_01011; 
		1465: oled_colour = 16'b00110_001110_01100; 
		1466: oled_colour = 16'b11001_101110_01001; 
		1467: oled_colour = 16'b11111_111100_00010; 
		1468: oled_colour = 16'b11111_111000_00011; 
		1469: oled_colour = 16'b11111_111000_00101; 
		1470: oled_colour = 16'b11101_110010_01010; 
		1471: oled_colour = 16'b10110_101010_01100; 
		1472: oled_colour = 16'b10000_011111_01101; 
		1473: oled_colour = 16'b01001_010011_01110; 
		1474: oled_colour = 16'b00100_001100_01101; 
		1475: oled_colour = 16'b00010_001010_01100; 
		1476: oled_colour = 16'b00011_001101_01101; 
		1477: oled_colour = 16'b00100_001110_01110; 
		1478: oled_colour = 16'b00101_001111_01110; 
		1479: oled_colour = 16'b00101_010000_01110; 
		1480: oled_colour = 16'b00100_010000_01101; 
		1481: oled_colour = 16'b00110_010011_01111; 
		1482: oled_colour = 16'b01000_010101_10000; 
		1483: oled_colour = 16'b01000_010101_10000; 
		1484: oled_colour = 16'b00111_010011_01111; 
		1485: oled_colour = 16'b00110_010001_01110; 
		1486: oled_colour = 16'b00101_001111_01110; 
		1487: oled_colour = 16'b00101_001110_01110; 
		1488: oled_colour = 16'b00101_001110_01110; 
		1489: oled_colour = 16'b00110_010011_10000; 
		1490: oled_colour = 16'b01010_011010_10001; 
		1491: oled_colour = 16'b01100_011100_10010; 
		1492: oled_colour = 16'b01011_011011_10010; 
		1493: oled_colour = 16'b01001_011001_10000; 
		1494: oled_colour = 16'b01000_010101_01111; 
		1495: oled_colour = 16'b01000_010110_10000; 
		1496: oled_colour = 16'b00111_010011_10000; 
		1497: oled_colour = 16'b00110_010001_01111; 
		1498: oled_colour = 16'b00100_001110_01101; 
		1499: oled_colour = 16'b00011_001010_01100; 
		1500: oled_colour = 16'b00010_000110_01011; 
		1501: oled_colour = 16'b00010_000101_01001; 
		1502: oled_colour = 16'b00011_000111_01010; 
		1503: oled_colour = 16'b00101_001011_01100; 
		1504: oled_colour = 16'b00011_000110_01010; 
		1505: oled_colour = 16'b00010_000101_01010; 
		1506: oled_colour = 16'b00011_000101_01001; 
		1507: oled_colour = 16'b00011_000101_01001; 
		1508: oled_colour = 16'b00011_000101_01001; 
		1509: oled_colour = 16'b00011_000101_01001; 
		1510: oled_colour = 16'b00010_000101_01010; 
		1511: oled_colour = 16'b00010_000101_01010; 
		1512: oled_colour = 16'b00010_000101_01010; 
		1513: oled_colour = 16'b00010_000101_01010; 
		1514: oled_colour = 16'b00011_000101_01010; 
		1515: oled_colour = 16'b00011_000101_01001; 
		1516: oled_colour = 16'b00011_000101_01001; 
		1517: oled_colour = 16'b00011_000101_01001; 
		1518: oled_colour = 16'b00011_000101_01001; 
		1519: oled_colour = 16'b00010_000101_01010; 
		1520: oled_colour = 16'b00010_000101_01010; 
		1521: oled_colour = 16'b00010_000110_01010; 
		1522: oled_colour = 16'b00010_000101_01001; 
		1523: oled_colour = 16'b00011_000111_01010; 
		1524: oled_colour = 16'b00110_001011_01000; 
		1525: oled_colour = 16'b00100_001001_00101; 
		1526: oled_colour = 16'b01100_011010_01101; 
		1527: oled_colour = 16'b01101_011101_01101; 
		1528: oled_colour = 16'b01101_011011_01101; 
		1529: oled_colour = 16'b01101_011010_01101; 
		1530: oled_colour = 16'b01001_010011_01010; 
		1531: oled_colour = 16'b01010_010110_01011; 
		1532: oled_colour = 16'b10010_100011_01111; 
		1533: oled_colour = 16'b00101_001100_01000; 
		1534: oled_colour = 16'b01001_010100_01011; 
		1535: oled_colour = 16'b10010_100011_01111; 
		1536: oled_colour = 16'b01010_010101_01001; 
		1537: oled_colour = 16'b01100_011000_01010; 
		1538: oled_colour = 16'b01111_011101_01011; 
		1539: oled_colour = 16'b00110_001010_01010; 
		1540: oled_colour = 16'b00001_000100_01011; 
		1541: oled_colour = 16'b00011_000110_01011; 
		1542: oled_colour = 16'b00010_000111_01011; 
		1543: oled_colour = 16'b00010_000111_01011; 
		1544: oled_colour = 16'b00010_000111_01011; 
		1545: oled_colour = 16'b00010_000110_01011; 
		1546: oled_colour = 16'b00010_000110_01011; 
		1547: oled_colour = 16'b00010_000110_01011; 
		1548: oled_colour = 16'b00010_000101_01011; 
		1549: oled_colour = 16'b00010_000101_01011; 
		1550: oled_colour = 16'b00010_000101_01011; 
		1551: oled_colour = 16'b00010_000101_01011; 
		1552: oled_colour = 16'b00010_000110_01011; 
		1553: oled_colour = 16'b00010_000110_01010; 
		1554: oled_colour = 16'b00010_000110_01011; 
		1555: oled_colour = 16'b00010_000110_01011; 
		1556: oled_colour = 16'b00011_000110_01011; 
		1557: oled_colour = 16'b00010_000110_01011; 
		1558: oled_colour = 16'b00010_000110_01011; 
		1559: oled_colour = 16'b00010_000110_01011; 
		1560: oled_colour = 16'b00010_000101_01011; 
		1561: oled_colour = 16'b00001_000110_01101; 
		1562: oled_colour = 16'b01001_010110_01110; 
		1563: oled_colour = 16'b11110_110111_00111; 
		1564: oled_colour = 16'b11111_111010_00011; 
		1565: oled_colour = 16'b11111_110110_00110; 
		1566: oled_colour = 16'b11101_110100_01001; 
		1567: oled_colour = 16'b11101_110011_01010; 
		1568: oled_colour = 16'b11010_101110_01110; 
		1569: oled_colour = 16'b10100_100100_10010; 
		1570: oled_colour = 16'b01110_011110_10010; 
		1571: oled_colour = 16'b01100_011101_10010; 
		1572: oled_colour = 16'b01101_011101_10010; 
		1573: oled_colour = 16'b01101_011110_10010; 
		1574: oled_colour = 16'b01100_011100_10010; 
		1575: oled_colour = 16'b01010_011001_10001; 
		1576: oled_colour = 16'b01000_010111_10000; 
		1577: oled_colour = 16'b00110_010100_01111; 
		1578: oled_colour = 16'b00101_010000_01110; 
		1579: oled_colour = 16'b00100_001110_01110; 
		1580: oled_colour = 16'b00100_001101_01110; 
		1581: oled_colour = 16'b00100_001101_01101; 
		1582: oled_colour = 16'b00011_001100_01101; 
		1583: oled_colour = 16'b00011_001001_01100; 
		1584: oled_colour = 16'b00010_001000_01100; 
		1585: oled_colour = 16'b00010_001010_01101; 
		1586: oled_colour = 16'b00100_001110_01110; 
		1587: oled_colour = 16'b00101_001110_01110; 
		1588: oled_colour = 16'b00111_010100_10000; 
		1589: oled_colour = 16'b01000_010111_10000; 
		1590: oled_colour = 16'b00110_010000_01101; 
		1591: oled_colour = 16'b00111_010010_01111; 
		1592: oled_colour = 16'b00111_010011_01111; 
		1593: oled_colour = 16'b01000_010011_10000; 
		1594: oled_colour = 16'b00101_010000_01101; 
		1595: oled_colour = 16'b00010_001010_01100; 
		1596: oled_colour = 16'b00010_000111_01100; 
		1597: oled_colour = 16'b00001_000100_01010; 
		1598: oled_colour = 16'b00110_001111_01101; 
		1599: oled_colour = 16'b00110_001111_01110; 
		1600: oled_colour = 16'b00010_000100_01010; 
		1601: oled_colour = 16'b00010_000110_01011; 
		1602: oled_colour = 16'b00010_000110_01011; 
		1603: oled_colour = 16'b00010_000101_01010; 
		1604: oled_colour = 16'b00010_000101_01010; 
		1605: oled_colour = 16'b00010_000101_01010; 
		1606: oled_colour = 16'b00010_000101_01010; 
		1607: oled_colour = 16'b00010_000101_01010; 
		1608: oled_colour = 16'b00010_000101_01011; 
		1609: oled_colour = 16'b00010_000101_01011; 
		1610: oled_colour = 16'b00010_000110_01011; 
		1611: oled_colour = 16'b00010_000110_01011; 
		1612: oled_colour = 16'b00010_000110_01010; 
		1613: oled_colour = 16'b00010_000101_01010; 
		1614: oled_colour = 16'b00010_000101_01010; 
		1615: oled_colour = 16'b00010_000101_01011; 
		1616: oled_colour = 16'b00010_000110_01011; 
		1617: oled_colour = 16'b00010_000110_01011; 
		1618: oled_colour = 16'b00010_000100_01010; 
		1619: oled_colour = 16'b00100_001001_01011; 
		1620: oled_colour = 16'b00111_001111_01001; 
		1621: oled_colour = 16'b00101_001010_00110; 
		1622: oled_colour = 16'b00111_010010_01011; 
		1623: oled_colour = 16'b00110_001111_01001; 
		1624: oled_colour = 16'b01000_010010_01010; 
		1625: oled_colour = 16'b01001_010100_01010; 
		1626: oled_colour = 16'b01001_010101_01011; 
		1627: oled_colour = 16'b01001_010100_01010; 
		1628: oled_colour = 16'b01110_011100_01101; 
		1629: oled_colour = 16'b00111_010000_01010; 
		1630: oled_colour = 16'b00111_010000_01001; 
		1631: oled_colour = 16'b01111_011111_01110; 
		1632: oled_colour = 16'b01011_010111_01010; 
		1633: oled_colour = 16'b01011_010110_01010; 
		1634: oled_colour = 16'b01110_011011_01010; 
		1635: oled_colour = 16'b01110_011000_01011; 
		1636: oled_colour = 16'b00001_000100_01010; 
		1637: oled_colour = 16'b00011_000110_01011; 
		1638: oled_colour = 16'b00010_000110_01011; 
		1639: oled_colour = 16'b00010_000110_01011; 
		1640: oled_colour = 16'b00010_000101_01011; 
		1641: oled_colour = 16'b00010_000101_01011; 
		1642: oled_colour = 16'b00011_000101_01011; 
		1643: oled_colour = 16'b00011_000110_01011; 
		1644: oled_colour = 16'b00011_000110_01011; 
		1645: oled_colour = 16'b00010_000110_01011; 
		1646: oled_colour = 16'b00010_000101_01011; 
		1647: oled_colour = 16'b00011_000101_01011; 
		1648: oled_colour = 16'b00010_000101_01011; 
		1649: oled_colour = 16'b00010_000101_01011; 
		1650: oled_colour = 16'b00010_000101_01011; 
		1651: oled_colour = 16'b00010_000101_01011; 
		1652: oled_colour = 16'b00010_000101_01011; 
		1653: oled_colour = 16'b00010_000101_01011; 
		1654: oled_colour = 16'b00010_000101_01011; 
		1655: oled_colour = 16'b00010_000101_01011; 
		1656: oled_colour = 16'b00010_000101_01011; 
		1657: oled_colour = 16'b00011_000110_01011; 
		1658: oled_colour = 16'b00010_001000_01100; 
		1659: oled_colour = 16'b01011_011010_01101; 
		1660: oled_colour = 16'b11011_110010_01001; 
		1661: oled_colour = 16'b11111_111010_00100; 
		1662: oled_colour = 16'b11111_111101_00010; 
		1663: oled_colour = 16'b11111_111100_00011; 
		1664: oled_colour = 16'b11111_111000_00111; 
		1665: oled_colour = 16'b11010_101101_01101; 
		1666: oled_colour = 16'b10000_100001_01101; 
		1667: oled_colour = 16'b01011_011010_10000; 
		1668: oled_colour = 16'b01001_010110_10000; 
		1669: oled_colour = 16'b01001_010110_10000; 
		1670: oled_colour = 16'b01000_010110_10000; 
		1671: oled_colour = 16'b01000_010110_10000; 
		1672: oled_colour = 16'b01001_010110_10000; 
		1673: oled_colour = 16'b01000_010101_10000; 
		1674: oled_colour = 16'b00111_010100_01111; 
		1675: oled_colour = 16'b00110_010010_01111; 
		1676: oled_colour = 16'b00101_010001_01110; 
		1677: oled_colour = 16'b00101_010000_01110; 
		1678: oled_colour = 16'b00100_001111_01110; 
		1679: oled_colour = 16'b00011_001101_01101; 
		1680: oled_colour = 16'b00010_001011_01101; 
		1681: oled_colour = 16'b00010_001001_01101; 
		1682: oled_colour = 16'b00010_000110_01100; 
		1683: oled_colour = 16'b00010_000101_01011; 
		1684: oled_colour = 16'b00100_001010_01101; 
		1685: oled_colour = 16'b00100_010000_01100; 
		1686: oled_colour = 16'b00011_001100_01100; 
		1687: oled_colour = 16'b00101_001111_01111; 
		1688: oled_colour = 16'b00101_001111_01111; 
		1689: oled_colour = 16'b00110_010001_10000; 
		1690: oled_colour = 16'b00110_010001_10000; 
		1691: oled_colour = 16'b00100_001100_01110; 
		1692: oled_colour = 16'b00100_001011_01101; 
		1693: oled_colour = 16'b00011_001001_01100; 
		1694: oled_colour = 16'b00100_001011_01011; 
		1695: oled_colour = 16'b00110_010010_01110; 
		1696: oled_colour = 16'b00010_000101_01011; 
		1697: oled_colour = 16'b00010_000110_01011; 
		1698: oled_colour = 16'b00010_000110_01011; 
		1699: oled_colour = 16'b00010_000110_01011; 
		1700: oled_colour = 16'b00010_000110_01011; 
		1701: oled_colour = 16'b00010_000110_01011; 
		1702: oled_colour = 16'b00010_000110_01011; 
		1703: oled_colour = 16'b00010_000110_01011; 
		1704: oled_colour = 16'b00010_000110_01011; 
		1705: oled_colour = 16'b00010_000110_01011; 
		1706: oled_colour = 16'b00010_000110_01011; 
		1707: oled_colour = 16'b00010_000110_01011; 
		1708: oled_colour = 16'b00010_000110_01011; 
		1709: oled_colour = 16'b00010_000110_01011; 
		1710: oled_colour = 16'b00010_000110_01011; 
		1711: oled_colour = 16'b00010_000110_01011; 
		1712: oled_colour = 16'b00010_000110_01011; 
		1713: oled_colour = 16'b00010_000110_01011; 
		1714: oled_colour = 16'b00010_000100_01010; 
		1715: oled_colour = 16'b00110_001101_01101; 
		1716: oled_colour = 16'b00100_001000_00100; 
		1717: oled_colour = 16'b00010_000101_00100; 
		1718: oled_colour = 16'b01100_011011_01101; 
		1719: oled_colour = 16'b01110_011110_01101; 
		1720: oled_colour = 16'b01110_011101_01101; 
		1721: oled_colour = 16'b01101_011011_01101; 
		1722: oled_colour = 16'b01010_010111_01011; 
		1723: oled_colour = 16'b00110_010000_01001; 
		1724: oled_colour = 16'b10000_100001_01111; 
		1725: oled_colour = 16'b01000_010010_01001; 
		1726: oled_colour = 16'b00101_001110_01001; 
		1727: oled_colour = 16'b01111_011111_01110; 
		1728: oled_colour = 16'b01110_011011_01010; 
		1729: oled_colour = 16'b01010_010101_01010; 
		1730: oled_colour = 16'b01100_011000_01010; 
		1731: oled_colour = 16'b10001_100000_01011; 
		1732: oled_colour = 16'b01000_001111_01010; 
		1733: oled_colour = 16'b00001_000011_01011; 
		1734: oled_colour = 16'b00010_000101_01011; 
		1735: oled_colour = 16'b00010_000100_01010; 
		1736: oled_colour = 16'b00001_000101_01011; 
		1737: oled_colour = 16'b00010_000110_01011; 
		1738: oled_colour = 16'b00001_000101_01011; 
		1739: oled_colour = 16'b00001_000110_01100; 
		1740: oled_colour = 16'b00010_001001_01100; 
		1741: oled_colour = 16'b00010_001010_01100; 
		1742: oled_colour = 16'b00010_000111_01100; 
		1743: oled_colour = 16'b00001_000110_01011; 
		1744: oled_colour = 16'b00010_000111_01100; 
		1745: oled_colour = 16'b00010_001000_01100; 
		1746: oled_colour = 16'b00010_001000_01100; 
		1747: oled_colour = 16'b00010_001001_01100; 
		1748: oled_colour = 16'b00010_001010_01100; 
		1749: oled_colour = 16'b00010_001001_01100; 
		1750: oled_colour = 16'b00010_001010_01100; 
		1751: oled_colour = 16'b00010_001010_01100; 
		1752: oled_colour = 16'b00010_001001_01100; 
		1753: oled_colour = 16'b00010_001000_01011; 
		1754: oled_colour = 16'b00010_001000_01100; 
		1755: oled_colour = 16'b00001_001000_01100; 
		1756: oled_colour = 16'b00011_001101_01110; 
		1757: oled_colour = 16'b01011_011001_01110; 
		1758: oled_colour = 16'b10010_100011_01011; 
		1759: oled_colour = 16'b10011_100110_01010; 
		1760: oled_colour = 16'b01111_011111_01011; 
		1761: oled_colour = 16'b00110_010001_01101; 
		1762: oled_colour = 16'b00001_001000_01100; 
		1763: oled_colour = 16'b00001_001001_01100; 
		1764: oled_colour = 16'b00010_001001_01100; 
		1765: oled_colour = 16'b00010_001001_01100; 
		1766: oled_colour = 16'b00010_001000_01100; 
		1767: oled_colour = 16'b00010_000110_01011; 
		1768: oled_colour = 16'b00010_000110_01011; 
		1769: oled_colour = 16'b00010_000110_01011; 
		1770: oled_colour = 16'b00010_000110_01011; 
		1771: oled_colour = 16'b00010_000101_01011; 
		1772: oled_colour = 16'b00010_000101_01011; 
		1773: oled_colour = 16'b00010_000101_01011; 
		1774: oled_colour = 16'b00010_000101_01011; 
		1775: oled_colour = 16'b00010_000110_01011; 
		1776: oled_colour = 16'b00010_000111_01100; 
		1777: oled_colour = 16'b00010_001000_01100; 
		1778: oled_colour = 16'b00011_001001_01100; 
		1779: oled_colour = 16'b00010_000110_01011; 
		1780: oled_colour = 16'b00110_010000_10000; 
		1781: oled_colour = 16'b00100_010001_01011; 
		1782: oled_colour = 16'b00010_001011_00111; 
		1783: oled_colour = 16'b00011_001101_01001; 
		1784: oled_colour = 16'b00011_001110_01001; 
		1785: oled_colour = 16'b00100_001111_01001; 
		1786: oled_colour = 16'b00101_010001_01011; 
		1787: oled_colour = 16'b00100_010000_01010; 
		1788: oled_colour = 16'b00100_001111_01010; 
		1789: oled_colour = 16'b00011_001110_01001; 
		1790: oled_colour = 16'b00011_001110_01001; 
		1791: oled_colour = 16'b00011_001011_01011; 
		1792: oled_colour = 16'b00010_000100_01011; 
		1793: oled_colour = 16'b00010_000110_01011; 
		1794: oled_colour = 16'b00010_000110_01011; 
		1795: oled_colour = 16'b00010_000110_01011; 
		1796: oled_colour = 16'b00010_000110_01011; 
		1797: oled_colour = 16'b00010_000110_01011; 
		1798: oled_colour = 16'b00010_000110_01011; 
		1799: oled_colour = 16'b00010_000110_01011; 
		1800: oled_colour = 16'b00010_000110_01011; 
		1801: oled_colour = 16'b00010_000110_01011; 
		1802: oled_colour = 16'b00010_000110_01011; 
		1803: oled_colour = 16'b00010_000110_01011; 
		1804: oled_colour = 16'b00010_000110_01011; 
		1805: oled_colour = 16'b00010_000110_01011; 
		1806: oled_colour = 16'b00010_000110_01011; 
		1807: oled_colour = 16'b00010_000110_01011; 
		1808: oled_colour = 16'b00010_000110_01011; 
		1809: oled_colour = 16'b00010_000110_01011; 
		1810: oled_colour = 16'b00010_000101_01011; 
		1811: oled_colour = 16'b00111_001110_01100; 
		1812: oled_colour = 16'b00100_000111_00100; 
		1813: oled_colour = 16'b00011_000110_00100; 
		1814: oled_colour = 16'b00111_010001_01010; 
		1815: oled_colour = 16'b01001_010100_01010; 
		1816: oled_colour = 16'b01010_010110_01011; 
		1817: oled_colour = 16'b01011_011000_01011; 
		1818: oled_colour = 16'b01100_011010_01100; 
		1819: oled_colour = 16'b01010_010101_01011; 
		1820: oled_colour = 16'b01110_011110_01110; 
		1821: oled_colour = 16'b01001_010011_01010; 
		1822: oled_colour = 16'b00101_001100_01000; 
		1823: oled_colour = 16'b01111_011110_01110; 
		1824: oled_colour = 16'b01111_011101_01010; 
		1825: oled_colour = 16'b01011_010111_01010; 
		1826: oled_colour = 16'b01100_010111_01010; 
		1827: oled_colour = 16'b01110_011011_01010; 
		1828: oled_colour = 16'b10000_011110_01010; 
		1829: oled_colour = 16'b00011_000111_01011; 
		1830: oled_colour = 16'b00011_001001_01100; 
		1831: oled_colour = 16'b00101_001110_01110; 
		1832: oled_colour = 16'b01000_010100_10000; 
		1833: oled_colour = 16'b01001_010111_10000; 
		1834: oled_colour = 16'b01001_010110_10000; 
		1835: oled_colour = 16'b01010_010110_10000; 
		1836: oled_colour = 16'b01010_010111_10000; 
		1837: oled_colour = 16'b01010_011001_10000; 
		1838: oled_colour = 16'b01011_011001_10000; 
		1839: oled_colour = 16'b01100_011011_10000; 
		1840: oled_colour = 16'b01100_011011_10000; 
		1841: oled_colour = 16'b01100_011011_10001; 
		1842: oled_colour = 16'b01100_011100_10001; 
		1843: oled_colour = 16'b01100_011011_10001; 
		1844: oled_colour = 16'b01100_011100_10001; 
		1845: oled_colour = 16'b01100_011100_10001; 
		1846: oled_colour = 16'b01100_011011_10001; 
		1847: oled_colour = 16'b01011_011010_10000; 
		1848: oled_colour = 16'b01011_011011_10001; 
		1849: oled_colour = 16'b01011_011011_10001; 
		1850: oled_colour = 16'b01011_011010_10001; 
		1851: oled_colour = 16'b01011_011001_10001; 
		1852: oled_colour = 16'b01001_010110_10000; 
		1853: oled_colour = 16'b01000_010110_10000; 
		1854: oled_colour = 16'b01000_010101_10000; 
		1855: oled_colour = 16'b01000_010100_10000; 
		1856: oled_colour = 16'b00111_010101_10000; 
		1857: oled_colour = 16'b01000_010110_10000; 
		1858: oled_colour = 16'b01010_011000_10000; 
		1859: oled_colour = 16'b01001_010111_10001; 
		1860: oled_colour = 16'b01000_010110_10000; 
		1861: oled_colour = 16'b00110_010011_01111; 
		1862: oled_colour = 16'b00011_001110_01101; 
		1863: oled_colour = 16'b00010_001001_01100; 
		1864: oled_colour = 16'b00010_000110_01011; 
		1865: oled_colour = 16'b00010_000101_01011; 
		1866: oled_colour = 16'b00010_000101_01011; 
		1867: oled_colour = 16'b00010_000101_01011; 
		1868: oled_colour = 16'b00010_000101_01011; 
		1869: oled_colour = 16'b00010_000101_01011; 
		1870: oled_colour = 16'b00010_000101_01011; 
		1871: oled_colour = 16'b00010_000101_01011; 
		1872: oled_colour = 16'b00010_000101_01011; 
		1873: oled_colour = 16'b00010_000101_01011; 
		1874: oled_colour = 16'b00010_000101_01011; 
		1875: oled_colour = 16'b00010_000100_01010; 
		1876: oled_colour = 16'b00101_001111_01110; 
		1877: oled_colour = 16'b00011_001111_01001; 
		1878: oled_colour = 16'b00001_001001_00110; 
		1879: oled_colour = 16'b00001_001001_00110; 
		1880: oled_colour = 16'b00001_001001_00110; 
		1881: oled_colour = 16'b00001_001001_00110; 
		1882: oled_colour = 16'b00001_001001_00101; 
		1883: oled_colour = 16'b00001_001001_00110; 
		1884: oled_colour = 16'b00001_001001_00110; 
		1885: oled_colour = 16'b00001_001001_00110; 
		1886: oled_colour = 16'b00010_001011_00110; 
		1887: oled_colour = 16'b00100_010001_01100; 
		1888: oled_colour = 16'b00011_001001_01100; 
		1889: oled_colour = 16'b00010_000100_01010; 
		1890: oled_colour = 16'b00010_000100_01010; 
		1891: oled_colour = 16'b00010_000101_01010; 
		1892: oled_colour = 16'b00010_000110_01011; 
		1893: oled_colour = 16'b00010_000101_01011; 
		1894: oled_colour = 16'b00010_000101_01011; 
		1895: oled_colour = 16'b00010_000110_01011; 
		1896: oled_colour = 16'b00010_000101_01011; 
		1897: oled_colour = 16'b00010_000101_01011; 
		1898: oled_colour = 16'b00010_000101_01011; 
		1899: oled_colour = 16'b00010_000101_01011; 
		1900: oled_colour = 16'b00010_000101_01011; 
		1901: oled_colour = 16'b00010_000101_01011; 
		1902: oled_colour = 16'b00010_000110_01011; 
		1903: oled_colour = 16'b00010_000101_01011; 
		1904: oled_colour = 16'b00010_000110_01011; 
		1905: oled_colour = 16'b00010_000101_01011; 
		1906: oled_colour = 16'b00011_000111_01011; 
		1907: oled_colour = 16'b00110_001101_01010; 
		1908: oled_colour = 16'b00011_000101_00010; 
		1909: oled_colour = 16'b00010_000011_00011; 
		1910: oled_colour = 16'b01000_010010_01001; 
		1911: oled_colour = 16'b01110_011110_01110; 
		1912: oled_colour = 16'b01101_011011_01101; 
		1913: oled_colour = 16'b01100_011010_01100; 
		1914: oled_colour = 16'b01011_011000_01100; 
		1915: oled_colour = 16'b00101_001110_01000; 
		1916: oled_colour = 16'b01111_011110_01110; 
		1917: oled_colour = 16'b01101_011010_01100; 
		1918: oled_colour = 16'b00011_001011_00111; 
		1919: oled_colour = 16'b01110_011100_01101; 
		1920: oled_colour = 16'b10100_100001_01011; 
		1921: oled_colour = 16'b01101_011011_01010; 
		1922: oled_colour = 16'b01010_010101_01010; 
		1923: oled_colour = 16'b01100_011000_01010; 
		1924: oled_colour = 16'b10000_011101_01010; 
		1925: oled_colour = 16'b01010_010100_01011; 
		1926: oled_colour = 16'b00010_001011_01101; 
		1927: oled_colour = 16'b00111_010100_10000; 
		1928: oled_colour = 16'b01010_011000_10000; 
		1929: oled_colour = 16'b01011_011001_10001; 
		1930: oled_colour = 16'b01011_011010_10001; 
		1931: oled_colour = 16'b01100_011100_10001; 
		1932: oled_colour = 16'b01101_011100_10001; 
		1933: oled_colour = 16'b01110_011110_10010; 
		1934: oled_colour = 16'b01110_011111_10010; 
		1935: oled_colour = 16'b10001_100010_10010; 
		1936: oled_colour = 16'b10010_100100_10010; 
		1937: oled_colour = 16'b10011_100100_10010; 
		1938: oled_colour = 16'b10010_100010_10010; 
		1939: oled_colour = 16'b10000_100000_10010; 
		1940: oled_colour = 16'b01110_011110_10010; 
		1941: oled_colour = 16'b01101_011100_10001; 
		1942: oled_colour = 16'b01101_011100_10010; 
		1943: oled_colour = 16'b01110_011111_10010; 
		1944: oled_colour = 16'b01111_100000_10010; 
		1945: oled_colour = 16'b01110_011101_10001; 
		1946: oled_colour = 16'b01100_011100_10001; 
		1947: oled_colour = 16'b01011_011010_10001; 
		1948: oled_colour = 16'b01011_011010_10001; 
		1949: oled_colour = 16'b01011_011010_10000; 
		1950: oled_colour = 16'b01100_011100_10001; 
		1951: oled_colour = 16'b01100_011100_10001; 
		1952: oled_colour = 16'b01100_011011_10001; 
		1953: oled_colour = 16'b01011_011010_10001; 
		1954: oled_colour = 16'b01010_011000_10001; 
		1955: oled_colour = 16'b01001_010111_10001; 
		1956: oled_colour = 16'b00111_010100_10000; 
		1957: oled_colour = 16'b00101_010001_01110; 
		1958: oled_colour = 16'b00011_001100_01101; 
		1959: oled_colour = 16'b00010_001000_01100; 
		1960: oled_colour = 16'b00010_001000_01100; 
		1961: oled_colour = 16'b00010_000111_01100; 
		1962: oled_colour = 16'b00010_000111_01100; 
		1963: oled_colour = 16'b00010_000111_01100; 
		1964: oled_colour = 16'b00010_000111_01100; 
		1965: oled_colour = 16'b00010_000111_01100; 
		1966: oled_colour = 16'b00010_000111_01100; 
		1967: oled_colour = 16'b00010_000111_01100; 
		1968: oled_colour = 16'b00010_000111_01100; 
		1969: oled_colour = 16'b00010_000111_01100; 
		1970: oled_colour = 16'b00011_000111_01100; 
		1971: oled_colour = 16'b00010_000111_01100; 
		1972: oled_colour = 16'b00111_010011_01111; 
		1973: oled_colour = 16'b00010_001010_00110; 
		1974: oled_colour = 16'b00001_001001_00101; 
		1975: oled_colour = 16'b00001_001000_00101; 
		1976: oled_colour = 16'b00010_001001_00101; 
		1977: oled_colour = 16'b00010_001010_00110; 
		1978: oled_colour = 16'b00001_001001_00101; 
		1979: oled_colour = 16'b00001_001000_00101; 
		1980: oled_colour = 16'b00010_001000_00101; 
		1981: oled_colour = 16'b00001_001000_00101; 
		1982: oled_colour = 16'b00001_001000_00101; 
		1983: oled_colour = 16'b00011_001100_01000; 
		1984: oled_colour = 16'b00111_010110_01111; 
		1985: oled_colour = 16'b00101_010010_01110; 
		1986: oled_colour = 16'b00101_001101_01110; 
		1987: oled_colour = 16'b00011_001001_01101; 
		1988: oled_colour = 16'b00010_000110_01011; 
		1989: oled_colour = 16'b00010_000111_01100; 
		1990: oled_colour = 16'b00010_000111_01100; 
		1991: oled_colour = 16'b00010_000111_01100; 
		1992: oled_colour = 16'b00010_000111_01100; 
		1993: oled_colour = 16'b00010_000111_01100; 
		1994: oled_colour = 16'b00010_000111_01100; 
		1995: oled_colour = 16'b00010_000111_01100; 
		1996: oled_colour = 16'b00010_000111_01100; 
		1997: oled_colour = 16'b00010_000111_01100; 
		1998: oled_colour = 16'b00010_000111_01100; 
		1999: oled_colour = 16'b00010_000111_01100; 
		2000: oled_colour = 16'b00011_000111_01100; 
		2001: oled_colour = 16'b00010_000110_01011; 
		2002: oled_colour = 16'b00100_001010_01101; 
		2003: oled_colour = 16'b00110_001011_01000; 
		2004: oled_colour = 16'b00010_000100_00010; 
		2005: oled_colour = 16'b00010_000100_00011; 
		2006: oled_colour = 16'b00110_001101_01000; 
		2007: oled_colour = 16'b01000_010011_01010; 
		2008: oled_colour = 16'b01001_010100_01010; 
		2009: oled_colour = 16'b01011_011000_01011; 
		2010: oled_colour = 16'b01101_011100_01100; 
		2011: oled_colour = 16'b01101_011101_01101; 
		2012: oled_colour = 16'b01100_011001_01100; 
		2013: oled_colour = 16'b01110_011101_01101; 
		2014: oled_colour = 16'b00101_001101_01000; 
		2015: oled_colour = 16'b01000_010011_01010; 
		2016: oled_colour = 16'b01101_011000_01001; 
		2017: oled_colour = 16'b01110_011100_01010; 
		2018: oled_colour = 16'b01001_010100_01010; 
		2019: oled_colour = 16'b01011_010110_01010; 
		2020: oled_colour = 16'b01101_011010_01010; 
		2021: oled_colour = 16'b10000_011101_01011; 
		2022: oled_colour = 16'b00110_010000_01100; 
		2023: oled_colour = 16'b00001_001011_01101; 
		2024: oled_colour = 16'b00010_001101_01101; 
		2025: oled_colour = 16'b00010_001100_01101; 
		2026: oled_colour = 16'b00011_001110_01101; 
		2027: oled_colour = 16'b00100_010000_01110; 
		2028: oled_colour = 16'b00101_010001_01110; 
		2029: oled_colour = 16'b00110_010010_01111; 
		2030: oled_colour = 16'b00111_010101_10000; 
		2031: oled_colour = 16'b01011_011010_10001; 
		2032: oled_colour = 16'b01111_011111_10010; 
		2033: oled_colour = 16'b10001_100010_10010; 
		2034: oled_colour = 16'b10010_100010_10010; 
		2035: oled_colour = 16'b10001_100010_10010; 
		2036: oled_colour = 16'b10000_100001_10010; 
		2037: oled_colour = 16'b01110_011110_10010; 
		2038: oled_colour = 16'b01110_011101_10010; 
		2039: oled_colour = 16'b01101_011100_10001; 
		2040: oled_colour = 16'b01100_011011_10001; 
		2041: oled_colour = 16'b01011_011010_10000; 
		2042: oled_colour = 16'b01001_011000_10000; 
		2043: oled_colour = 16'b01001_010110_10000; 
		2044: oled_colour = 16'b00111_010100_01111; 
		2045: oled_colour = 16'b00101_010001_01110; 
		2046: oled_colour = 16'b00011_001110_01101; 
		2047: oled_colour = 16'b00010_001101_01101; 
		2048: oled_colour = 16'b00010_001101_01101; 
		2049: oled_colour = 16'b00010_001011_01101; 
		2050: oled_colour = 16'b00010_001001_01101; 
		2051: oled_colour = 16'b00010_001010_01101; 
		2052: oled_colour = 16'b00010_001011_01101; 
		2053: oled_colour = 16'b00010_001011_01101; 
		2054: oled_colour = 16'b00010_001001_01101; 
		2055: oled_colour = 16'b00010_001001_01101; 
		2056: oled_colour = 16'b00010_001001_01101; 
		2057: oled_colour = 16'b00010_001001_01101; 
		2058: oled_colour = 16'b00010_001001_01101; 
		2059: oled_colour = 16'b00010_001001_01101; 
		2060: oled_colour = 16'b00010_001001_01101; 
		2061: oled_colour = 16'b00010_001001_01101; 
		2062: oled_colour = 16'b00010_001001_01101; 
		2063: oled_colour = 16'b00010_001001_01101; 
		2064: oled_colour = 16'b00010_001001_01101; 
		2065: oled_colour = 16'b00010_001001_01101; 
		2066: oled_colour = 16'b00010_001001_01101; 
		2067: oled_colour = 16'b00011_001100_01110; 
		2068: oled_colour = 16'b01000_011001_10001; 
		2069: oled_colour = 16'b00011_001010_00110; 
		2070: oled_colour = 16'b00010_001001_00110; 
		2071: oled_colour = 16'b00010_001011_00111; 
		2072: oled_colour = 16'b00011_001100_00111; 
		2073: oled_colour = 16'b00011_001100_00111; 
		2074: oled_colour = 16'b00001_001001_00101; 
		2075: oled_colour = 16'b00001_000111_00101; 
		2076: oled_colour = 16'b00010_001010_00110; 
		2077: oled_colour = 16'b00011_001010_00110; 
		2078: oled_colour = 16'b00001_001000_00101; 
		2079: oled_colour = 16'b00010_001000_00101; 
		2080: oled_colour = 16'b00011_001010_00110; 
		2081: oled_colour = 16'b00010_001011_00110; 
		2082: oled_colour = 16'b00111_010110_01111; 
		2083: oled_colour = 16'b00100_001101_01111; 
		2084: oled_colour = 16'b00010_001001_01101; 
		2085: oled_colour = 16'b00010_001010_01101; 
		2086: oled_colour = 16'b00010_001001_01101; 
		2087: oled_colour = 16'b00010_001001_01101; 
		2088: oled_colour = 16'b00010_001010_01101; 
		2089: oled_colour = 16'b00010_001010_01101; 
		2090: oled_colour = 16'b00010_001010_01101; 
		2091: oled_colour = 16'b00010_001010_01101; 
		2092: oled_colour = 16'b00010_001001_01101; 
		2093: oled_colour = 16'b00010_001001_01101; 
		2094: oled_colour = 16'b00010_001001_01101; 
		2095: oled_colour = 16'b00010_001001_01101; 
		2096: oled_colour = 16'b00010_001001_01101; 
		2097: oled_colour = 16'b00001_001001_01101; 
		2098: oled_colour = 16'b00101_001110_01110; 
		2099: oled_colour = 16'b00101_001010_00110; 
		2100: oled_colour = 16'b00010_000100_00011; 
		2101: oled_colour = 16'b00010_000100_00010; 
		2102: oled_colour = 16'b00101_001011_00110; 
		2103: oled_colour = 16'b01111_011111_01111; 
		2104: oled_colour = 16'b01110_011101_01110; 
		2105: oled_colour = 16'b01101_011011_01101; 
		2106: oled_colour = 16'b01100_011001_01100; 
		2107: oled_colour = 16'b01000_010011_01010; 
		2108: oled_colour = 16'b01000_010011_01010; 
		2109: oled_colour = 16'b10101_101001_10001; 
		2110: oled_colour = 16'b00111_001111_01001; 
		2111: oled_colour = 16'b00110_001111_01001; 
		2112: oled_colour = 16'b00111_001111_01001; 
		2113: oled_colour = 16'b01010_010011_01010; 
		2114: oled_colour = 16'b00111_001111_01001; 
		2115: oled_colour = 16'b00111_001101_00111; 
		2116: oled_colour = 16'b01100_011000_01010; 
		2117: oled_colour = 16'b01101_011010_01010; 
		2118: oled_colour = 16'b10001_100000_01100; 
		2119: oled_colour = 16'b01101_011100_10001; 
		2120: oled_colour = 16'b01100_011100_10001; 
		2121: oled_colour = 16'b01101_011101_10001; 
		2122: oled_colour = 16'b01110_011101_10001; 
		2123: oled_colour = 16'b01110_011111_10010; 
		2124: oled_colour = 16'b01111_100000_10010; 
		2125: oled_colour = 16'b10000_100000_10010; 
		2126: oled_colour = 16'b10000_100001_10010; 
		2127: oled_colour = 16'b10001_100001_10010; 
		2128: oled_colour = 16'b10010_100011_10010; 
		2129: oled_colour = 16'b10010_100011_10010; 
		2130: oled_colour = 16'b10001_100001_10010; 
		2131: oled_colour = 16'b01111_011111_10001; 
		2132: oled_colour = 16'b01110_011101_10001; 
		2133: oled_colour = 16'b01101_011100_10001; 
		2134: oled_colour = 16'b01100_011011_10001; 
		2135: oled_colour = 16'b01011_011001_10000; 
		2136: oled_colour = 16'b01010_011000_10000; 
		2137: oled_colour = 16'b01010_011000_10000; 
		2138: oled_colour = 16'b01001_010111_10000; 
		2139: oled_colour = 16'b01001_010111_10000; 
		2140: oled_colour = 16'b01000_010101_10000; 
		2141: oled_colour = 16'b00110_010011_01111; 
		2142: oled_colour = 16'b00011_001101_01101; 
		2143: oled_colour = 16'b00010_001011_01101; 
		2144: oled_colour = 16'b00011_001100_01101; 
		2145: oled_colour = 16'b00010_001010_01101; 
		2146: oled_colour = 16'b00010_001001_01101; 
		2147: oled_colour = 16'b00010_001001_01101; 
		2148: oled_colour = 16'b00010_001001_01101; 
		2149: oled_colour = 16'b00010_001001_01101; 
		2150: oled_colour = 16'b00010_001001_01101; 
		2151: oled_colour = 16'b00010_001001_01101; 
		2152: oled_colour = 16'b00010_001001_01101; 
		2153: oled_colour = 16'b00010_001001_01101; 
		2154: oled_colour = 16'b00010_001001_01101; 
		2155: oled_colour = 16'b00010_001001_01101; 
		2156: oled_colour = 16'b00010_001001_01101; 
		2157: oled_colour = 16'b00010_001001_01101; 
		2158: oled_colour = 16'b00010_001001_01101; 
		2159: oled_colour = 16'b00010_001001_01101; 
		2160: oled_colour = 16'b00010_001001_01101; 
		2161: oled_colour = 16'b00010_001010_01101; 
		2162: oled_colour = 16'b00001_000111_01100; 
		2163: oled_colour = 16'b00110_010110_10001; 
		2164: oled_colour = 16'b00100_010000_01010; 
		2165: oled_colour = 16'b00010_001000_00110; 
		2166: oled_colour = 16'b00110_010001_01011; 
		2167: oled_colour = 16'b00100_001110_01001; 
		2168: oled_colour = 16'b00011_001110_01001; 
		2169: oled_colour = 16'b00100_001110_01001; 
		2170: oled_colour = 16'b00100_001110_01001; 
		2171: oled_colour = 16'b00011_001101_01000; 
		2172: oled_colour = 16'b00011_001110_01001; 
		2173: oled_colour = 16'b00011_001110_01001; 
		2174: oled_colour = 16'b00011_001110_01001; 
		2175: oled_colour = 16'b00011_001101_01000; 
		2176: oled_colour = 16'b00100_001110_01000; 
		2177: oled_colour = 16'b00100_010000_01010; 
		2178: oled_colour = 16'b00011_001100_01101; 
		2179: oled_colour = 16'b00010_001000_01101; 
		2180: oled_colour = 16'b00010_001010_01101; 
		2181: oled_colour = 16'b00010_001001_01101; 
		2182: oled_colour = 16'b00010_001001_01101; 
		2183: oled_colour = 16'b00010_001001_01101; 
		2184: oled_colour = 16'b00010_001001_01101; 
		2185: oled_colour = 16'b00010_001001_01101; 
		2186: oled_colour = 16'b00010_001001_01101; 
		2187: oled_colour = 16'b00010_001001_01101; 
		2188: oled_colour = 16'b00010_001001_01101; 
		2189: oled_colour = 16'b00010_001010_01101; 
		2190: oled_colour = 16'b00011_001100_01101; 
		2191: oled_colour = 16'b00100_001110_01101; 
		2192: oled_colour = 16'b00101_010010_01110; 
		2193: oled_colour = 16'b01000_010110_10000; 
		2194: oled_colour = 16'b01000_010100_01110; 
		2195: oled_colour = 16'b00011_000101_00011; 
		2196: oled_colour = 16'b00010_000100_00011; 
		2197: oled_colour = 16'b00011_000100_00010; 
		2198: oled_colour = 16'b00011_000111_00100; 
		2199: oled_colour = 16'b01001_010100_01011; 
		2200: oled_colour = 16'b01010_010110_01011; 
		2201: oled_colour = 16'b01011_011001_01100; 
		2202: oled_colour = 16'b01100_011010_01100; 
		2203: oled_colour = 16'b01101_011101_01101; 
		2204: oled_colour = 16'b01001_010100_01010; 
		2205: oled_colour = 16'b10010_100101_01111; 
		2206: oled_colour = 16'b01000_010011_01010; 
		2207: oled_colour = 16'b00101_001100_01000; 
		2208: oled_colour = 16'b11000_110000_10010; 
		2209: oled_colour = 16'b10011_100101_01111; 
		2210: oled_colour = 16'b01011_011000_01100; 
		2211: oled_colour = 16'b00110_001101_01000; 
		2212: oled_colour = 16'b01001_010100_01010; 
		2213: oled_colour = 16'b01011_011000_01010; 
		2214: oled_colour = 16'b01110_011011_01010; 
		2215: oled_colour = 16'b10101_100110_01111; 
		2216: oled_colour = 16'b10010_100011_10010; 
		2217: oled_colour = 16'b10010_100011_10010; 
		2218: oled_colour = 16'b10011_100101_10010; 
		2219: oled_colour = 16'b10010_100100_10010; 
		2220: oled_colour = 16'b10001_100010_10010; 
		2221: oled_colour = 16'b10000_100000_10001; 
		2222: oled_colour = 16'b01101_011100_10001; 
		2223: oled_colour = 16'b01101_011100_10010; 
		2224: oled_colour = 16'b01011_011011_10001; 
		2225: oled_colour = 16'b01011_011011_10001; 
		2226: oled_colour = 16'b01100_011100_10010; 
		2227: oled_colour = 16'b01000_010101_10000; 
		2228: oled_colour = 16'b00101_010010_01110; 
		2229: oled_colour = 16'b00101_010001_01110; 
		2230: oled_colour = 16'b00011_001111_01101; 
		2231: oled_colour = 16'b00010_001101_01101; 
		2232: oled_colour = 16'b00010_001100_01101; 
		2233: oled_colour = 16'b00010_001011_01101; 
		2234: oled_colour = 16'b00001_001011_01100; 
		2235: oled_colour = 16'b00001_001010_01100; 
		2236: oled_colour = 16'b00001_001001_01100; 
		2237: oled_colour = 16'b00001_001001_01100; 
		2238: oled_colour = 16'b00010_001001_01100; 
		2239: oled_colour = 16'b00010_001010_01101; 
		2240: oled_colour = 16'b00010_001001_01101; 
		2241: oled_colour = 16'b00010_001001_01101; 
		2242: oled_colour = 16'b00010_001001_01101; 
		2243: oled_colour = 16'b00010_001001_01101; 
		2244: oled_colour = 16'b00010_001001_01101; 
		2245: oled_colour = 16'b00010_001001_01101; 
		2246: oled_colour = 16'b00010_001001_01101; 
		2247: oled_colour = 16'b00010_001001_01101; 
		2248: oled_colour = 16'b00010_001001_01101; 
		2249: oled_colour = 16'b00010_001001_01101; 
		2250: oled_colour = 16'b00010_001001_01101; 
		2251: oled_colour = 16'b00010_001001_01101; 
		2252: oled_colour = 16'b00010_001001_01101; 
		2253: oled_colour = 16'b00010_001001_01101; 
		2254: oled_colour = 16'b00010_001001_01101; 
		2255: oled_colour = 16'b00010_001001_01101; 
		2256: oled_colour = 16'b00010_001001_01101; 
		2257: oled_colour = 16'b00010_001000_01101; 
		2258: oled_colour = 16'b00100_001110_01110; 
		2259: oled_colour = 16'b00110_010111_01111; 
		2260: oled_colour = 16'b00001_000110_00100; 
		2261: oled_colour = 16'b00100_001101_01000; 
		2262: oled_colour = 16'b01000_010100_01100; 
		2263: oled_colour = 16'b00010_001001_00110; 
		2264: oled_colour = 16'b00010_001010_00110; 
		2265: oled_colour = 16'b00011_001011_00111; 
		2266: oled_colour = 16'b00010_001010_00110; 
		2267: oled_colour = 16'b00010_001001_00101; 
		2268: oled_colour = 16'b00010_001001_00110; 
		2269: oled_colour = 16'b00010_001001_00110; 
		2270: oled_colour = 16'b00010_001010_00110; 
		2271: oled_colour = 16'b00100_001110_01000; 
		2272: oled_colour = 16'b00100_001100_00111; 
		2273: oled_colour = 16'b00101_010000_01100; 
		2274: oled_colour = 16'b00011_001010_01101; 
		2275: oled_colour = 16'b00010_001001_01101; 
		2276: oled_colour = 16'b00010_001001_01101; 
		2277: oled_colour = 16'b00010_001001_01101; 
		2278: oled_colour = 16'b00010_001001_01101; 
		2279: oled_colour = 16'b00010_001001_01101; 
		2280: oled_colour = 16'b00010_001001_01101; 
		2281: oled_colour = 16'b00010_001001_01101; 
		2282: oled_colour = 16'b00010_001001_01101; 
		2283: oled_colour = 16'b00010_001001_01101; 
		2284: oled_colour = 16'b00010_001001_01101; 
		2285: oled_colour = 16'b00011_001101_01110; 
		2286: oled_colour = 16'b01000_010101_10000; 
		2287: oled_colour = 16'b01110_011101_10010; 
		2288: oled_colour = 16'b10001_100010_10010; 
		2289: oled_colour = 16'b10011_100101_10011; 
		2290: oled_colour = 16'b01010_010011_01011; 
		2291: oled_colour = 16'b00010_000011_00010; 
		2292: oled_colour = 16'b00011_000101_00011; 
		2293: oled_colour = 16'b00011_000101_00010; 
		2294: oled_colour = 16'b00010_000100_00011; 
		2295: oled_colour = 16'b01011_011000_01100; 
		2296: oled_colour = 16'b01111_100000_01110; 
		2297: oled_colour = 16'b01110_011100_01101; 
		2298: oled_colour = 16'b01101_011100_01101; 
		2299: oled_colour = 16'b01011_011000_01100; 
		2300: oled_colour = 16'b00111_010001_01001; 
		2301: oled_colour = 16'b01111_100000_01110; 
		2302: oled_colour = 16'b01101_011100_01101; 
		2303: oled_colour = 16'b00100_001100_01000; 
		2304: oled_colour = 16'b11100_110110_10011; 
		2305: oled_colour = 16'b11110_111001_10100; 
		2306: oled_colour = 16'b11100_110110_10011; 
		2307: oled_colour = 16'b11000_101111_10010; 
		2308: oled_colour = 16'b01010_010110_01011; 
		2309: oled_colour = 16'b00111_010000_01010; 
		2310: oled_colour = 16'b01000_010011_01001; 
		2311: oled_colour = 16'b01110_011011_01010; 
		2312: oled_colour = 16'b10010_100010_10000; 
		2313: oled_colour = 16'b01111_011111_10010; 
		2314: oled_colour = 16'b01111_100000_10010; 
		2315: oled_colour = 16'b01110_011110_10010; 
		2316: oled_colour = 16'b01101_011100_10001; 
		2317: oled_colour = 16'b01101_011100_10001; 
		2318: oled_colour = 16'b01101_011101_10010; 
		2319: oled_colour = 16'b01110_011111_10010; 
		2320: oled_colour = 16'b10000_100001_10010; 
		2321: oled_colour = 16'b10000_100001_10010; 
		2322: oled_colour = 16'b10001_100010_10010; 
		2323: oled_colour = 16'b10010_100010_10010; 
		2324: oled_colour = 16'b10001_100010_10010; 
		2325: oled_colour = 16'b10000_100001_10010; 
		2326: oled_colour = 16'b01111_100000_10010; 
		2327: oled_colour = 16'b01111_011111_10010; 
		2328: oled_colour = 16'b01110_011110_10010; 
		2329: oled_colour = 16'b01101_011101_10010; 
		2330: oled_colour = 16'b01101_011101_10001; 
		2331: oled_colour = 16'b01100_011011_10001; 
		2332: oled_colour = 16'b01011_011010_10001; 
		2333: oled_colour = 16'b01010_011000_10000; 
		2334: oled_colour = 16'b01001_010111_10000; 
		2335: oled_colour = 16'b01000_010110_10000; 
		2336: oled_colour = 16'b00111_010011_01111; 
		2337: oled_colour = 16'b00100_001111_01101; 
		2338: oled_colour = 16'b00011_001101_01101; 
		2339: oled_colour = 16'b00010_001100_01101; 
		2340: oled_colour = 16'b00010_001011_01101; 
		2341: oled_colour = 16'b00010_001011_01101; 
		2342: oled_colour = 16'b00010_001011_01101; 
		2343: oled_colour = 16'b00010_001011_01101; 
		2344: oled_colour = 16'b00010_001011_01101; 
		2345: oled_colour = 16'b00010_001011_01101; 
		2346: oled_colour = 16'b00010_001011_01101; 
		2347: oled_colour = 16'b00010_001011_01101; 
		2348: oled_colour = 16'b00010_001011_01101; 
		2349: oled_colour = 16'b00010_001011_01101; 
		2350: oled_colour = 16'b00010_001011_01101; 
		2351: oled_colour = 16'b00010_001011_01101; 
		2352: oled_colour = 16'b00010_001011_01101; 
		2353: oled_colour = 16'b00010_001010_01101; 
		2354: oled_colour = 16'b00101_010011_01111; 
		2355: oled_colour = 16'b00100_010010_01011; 
		2356: oled_colour = 16'b00001_000101_00011; 
		2357: oled_colour = 16'b00101_001110_01000; 
		2358: oled_colour = 16'b01001_010110_01101; 
		2359: oled_colour = 16'b00010_001010_00110; 
		2360: oled_colour = 16'b00101_001111_01001; 
		2361: oled_colour = 16'b00101_001111_01001; 
		2362: oled_colour = 16'b00010_001001_00101; 
		2363: oled_colour = 16'b00001_000110_00100; 
		2364: oled_colour = 16'b00001_000110_00100; 
		2365: oled_colour = 16'b00011_001100_01000; 
		2366: oled_colour = 16'b00100_001100_00111; 
		2367: oled_colour = 16'b00101_001111_01001; 
		2368: oled_colour = 16'b00100_001101_01000; 
		2369: oled_colour = 16'b00111_010100_01101; 
		2370: oled_colour = 16'b00010_001011_01101; 
		2371: oled_colour = 16'b00010_001011_01101; 
		2372: oled_colour = 16'b00010_001011_01101; 
		2373: oled_colour = 16'b00010_001011_01101; 
		2374: oled_colour = 16'b00010_001011_01101; 
		2375: oled_colour = 16'b00010_001011_01101; 
		2376: oled_colour = 16'b00010_001011_01101; 
		2377: oled_colour = 16'b00010_001011_01101; 
		2378: oled_colour = 16'b00010_001011_01101; 
		2379: oled_colour = 16'b00010_001011_01101; 
		2380: oled_colour = 16'b00010_001011_01101; 
		2381: oled_colour = 16'b00011_001101_01101; 
		2382: oled_colour = 16'b00110_010010_01110; 
		2383: oled_colour = 16'b01000_010110_10000; 
		2384: oled_colour = 16'b01010_011001_10001; 
		2385: oled_colour = 16'b01100_011011_10001; 
		2386: oled_colour = 16'b00111_001110_01001; 
		2387: oled_colour = 16'b00010_000011_00010; 
		2388: oled_colour = 16'b00011_000101_00010; 
		2389: oled_colour = 16'b00011_000101_00010; 
		2390: oled_colour = 16'b00010_000011_00011; 
		2391: oled_colour = 16'b00111_010001_01001; 
		2392: oled_colour = 16'b01111_100000_01110; 
		2393: oled_colour = 16'b01110_011110_01110; 
		2394: oled_colour = 16'b01111_011111_01101; 
		2395: oled_colour = 16'b01110_011110_01110; 
		2396: oled_colour = 16'b01011_011000_01100; 
		2397: oled_colour = 16'b01011_011000_01100; 
		2398: oled_colour = 16'b10010_100011_01111; 
		2399: oled_colour = 16'b00101_001101_01000; 
		2400: oled_colour = 16'b01011_010111_01011; 
		2401: oled_colour = 16'b10010_100100_01111; 
		2402: oled_colour = 16'b11001_110000_10010; 
		2403: oled_colour = 16'b11011_110100_10011; 
		2404: oled_colour = 16'b01100_011000_01100; 
		2405: oled_colour = 16'b10000_100010_01111; 
		2406: oled_colour = 16'b01011_010111_01100; 
		2407: oled_colour = 16'b00110_001110_01001; 
		2408: oled_colour = 16'b01001_010011_01010; 
		2409: oled_colour = 16'b00110_010010_01110; 
		2410: oled_colour = 16'b00100_010000_01110; 
		2411: oled_colour = 16'b00101_010001_01110; 
		2412: oled_colour = 16'b00101_010001_01110; 
		2413: oled_colour = 16'b00101_010010_01110; 
		2414: oled_colour = 16'b00110_010011_01111; 
		2415: oled_colour = 16'b00110_010100_01111; 
		2416: oled_colour = 16'b01000_010110_10000; 
		2417: oled_colour = 16'b01000_010101_01111; 
		2418: oled_colour = 16'b01001_010111_10000; 
		2419: oled_colour = 16'b01011_011001_10000; 
		2420: oled_colour = 16'b01010_011001_10000; 
		2421: oled_colour = 16'b01010_011000_10000; 
		2422: oled_colour = 16'b01001_010111_10000; 
		2423: oled_colour = 16'b01000_010110_10000; 
		2424: oled_colour = 16'b01000_010110_10000; 
		2425: oled_colour = 16'b00111_010101_01111; 
		2426: oled_colour = 16'b01000_010110_01111; 
		2427: oled_colour = 16'b01001_011000_10000; 
		2428: oled_colour = 16'b01001_010111_10000; 
		2429: oled_colour = 16'b00111_010101_01111; 
		2430: oled_colour = 16'b00111_010100_01111; 
		2431: oled_colour = 16'b00110_010011_01110; 
		2432: oled_colour = 16'b00101_010001_01101; 
		2433: oled_colour = 16'b00100_001111_01101; 
		2434: oled_colour = 16'b00011_001110_01101; 
		2435: oled_colour = 16'b00010_001101_01101; 
		2436: oled_colour = 16'b00010_001100_01101; 
		2437: oled_colour = 16'b00010_001100_01101; 
		2438: oled_colour = 16'b00010_001101_01101; 
		2439: oled_colour = 16'b00010_001100_01101; 
		2440: oled_colour = 16'b00010_001100_01101; 
		2441: oled_colour = 16'b00010_001100_01101; 
		2442: oled_colour = 16'b00010_001100_01101; 
		2443: oled_colour = 16'b00010_001100_01101; 
		2444: oled_colour = 16'b00010_001100_01101; 
		2445: oled_colour = 16'b00010_001100_01101; 
		2446: oled_colour = 16'b00010_001100_01101; 
		2447: oled_colour = 16'b00010_001101_01101; 
		2448: oled_colour = 16'b00010_001100_01101; 
		2449: oled_colour = 16'b00010_001100_01101; 
		2450: oled_colour = 16'b00001_001001_01100; 
		2451: oled_colour = 16'b00101_010101_10001; 
		2452: oled_colour = 16'b00100_001111_01001; 
		2453: oled_colour = 16'b00010_001010_00110; 
		2454: oled_colour = 16'b00111_010011_01100; 
		2455: oled_colour = 16'b00101_010000_01010; 
		2456: oled_colour = 16'b00011_001101_01001; 
		2457: oled_colour = 16'b00011_001101_01001; 
		2458: oled_colour = 16'b00011_001101_01001; 
		2459: oled_colour = 16'b00010_001100_01000; 
		2460: oled_colour = 16'b00100_001110_01000; 
		2461: oled_colour = 16'b00011_001100_01000; 
		2462: oled_colour = 16'b00110_001111_01001; 
		2463: oled_colour = 16'b00100_001101_01001; 
		2464: oled_colour = 16'b00101_001111_01010; 
		2465: oled_colour = 16'b01000_011000_01111; 
		2466: oled_colour = 16'b00011_010000_01110; 
		2467: oled_colour = 16'b00010_001011_01100; 
		2468: oled_colour = 16'b00001_001011_01100; 
		2469: oled_colour = 16'b00010_001100_01101; 
		2470: oled_colour = 16'b00010_001100_01101; 
		2471: oled_colour = 16'b00010_001100_01101; 
		2472: oled_colour = 16'b00010_001100_01101; 
		2473: oled_colour = 16'b00010_001100_01101; 
		2474: oled_colour = 16'b00010_001100_01101; 
		2475: oled_colour = 16'b00010_001100_01101; 
		2476: oled_colour = 16'b00010_001100_01101; 
		2477: oled_colour = 16'b00010_001100_01101; 
		2478: oled_colour = 16'b00010_001101_01101; 
		2479: oled_colour = 16'b00010_001101_01101; 
		2480: oled_colour = 16'b00011_001110_01101; 
		2481: oled_colour = 16'b00111_010011_01110; 
		2482: oled_colour = 16'b00011_000110_00100; 
		2483: oled_colour = 16'b00010_000101_00011; 
		2484: oled_colour = 16'b00010_000110_00100; 
		2485: oled_colour = 16'b00011_000110_00100; 
		2486: oled_colour = 16'b00010_000100_00011; 
		2487: oled_colour = 16'b00110_001101_01000; 
		2488: oled_colour = 16'b01110_011110_01110; 
		2489: oled_colour = 16'b01100_011001_01100; 
		2490: oled_colour = 16'b01110_011100_01101; 
		2491: oled_colour = 16'b01110_011100_01101; 
		2492: oled_colour = 16'b01101_011011_01100; 
		2493: oled_colour = 16'b01000_010010_01001; 
		2494: oled_colour = 16'b01111_011110_01110; 
		2495: oled_colour = 16'b00111_010001_01001; 
		2496: oled_colour = 16'b00010_000100_00011; 
		2497: oled_colour = 16'b00001_000011_00011; 
		2498: oled_colour = 16'b00110_001110_01001; 
		2499: oled_colour = 16'b01011_011001_01100; 
		2500: oled_colour = 16'b01011_011000_01100; 
		2501: oled_colour = 16'b11011_110101_10011; 
		2502: oled_colour = 16'b11011_110101_10011; 
		2503: oled_colour = 16'b10100_101000_10000; 
		2504: oled_colour = 16'b01100_011001_01100; 
		2505: oled_colour = 16'b00110_010000_01011; 
		2506: oled_colour = 16'b00011_001101_01100; 
		2507: oled_colour = 16'b00010_001100_01101; 
		2508: oled_colour = 16'b00011_001101_01101; 
		2509: oled_colour = 16'b00011_001101_01101; 
		2510: oled_colour = 16'b00010_001101_01101; 
		2511: oled_colour = 16'b00010_001101_01101; 
		2512: oled_colour = 16'b00010_001100_01101; 
		2513: oled_colour = 16'b00010_001100_01101; 
		2514: oled_colour = 16'b00010_001100_01101; 
		2515: oled_colour = 16'b00010_001011_01101; 
		2516: oled_colour = 16'b00001_001100_01101; 
		2517: oled_colour = 16'b00010_001100_01101; 
		2518: oled_colour = 16'b00010_001100_01101; 
		2519: oled_colour = 16'b00010_001100_01101; 
		2520: oled_colour = 16'b00010_001100_01101; 
		2521: oled_colour = 16'b00010_001100_01101; 
		2522: oled_colour = 16'b00010_001100_01101; 
		2523: oled_colour = 16'b00010_001101_01101; 
		2524: oled_colour = 16'b00010_001101_01101; 
		2525: oled_colour = 16'b00010_001101_01101; 
		2526: oled_colour = 16'b00011_001101_01101; 
		2527: oled_colour = 16'b00011_001101_01101; 
		2528: oled_colour = 16'b00011_001110_01101; 
		2529: oled_colour = 16'b00011_001110_01101; 
		2530: oled_colour = 16'b00010_001101_01101; 
		2531: oled_colour = 16'b00010_001100_01101; 
		2532: oled_colour = 16'b00010_001100_01101; 
		2533: oled_colour = 16'b00010_001100_01101; 
		2534: oled_colour = 16'b00010_001100_01101; 
		2535: oled_colour = 16'b00010_001100_01101; 
		2536: oled_colour = 16'b00010_001100_01101; 
		2537: oled_colour = 16'b00010_001100_01101; 
		2538: oled_colour = 16'b00010_001100_01101; 
		2539: oled_colour = 16'b00010_001100_01101; 
		2540: oled_colour = 16'b00010_001100_01101; 
		2541: oled_colour = 16'b00010_001101_01101; 
		2542: oled_colour = 16'b00011_001110_01110; 
		2543: oled_colour = 16'b00010_001100_01100; 
		2544: oled_colour = 16'b00010_001100_01101; 
		2545: oled_colour = 16'b00011_001110_01110; 
		2546: oled_colour = 16'b00100_010010_01111; 
		2547: oled_colour = 16'b01000_011010_10010; 
		2548: oled_colour = 16'b00100_001111_01010; 
		2549: oled_colour = 16'b00001_001001_00101; 
		2550: oled_colour = 16'b00001_001001_00110; 
		2551: oled_colour = 16'b00010_001010_00110; 
		2552: oled_colour = 16'b00010_001010_00111; 
		2553: oled_colour = 16'b00010_001010_00110; 
		2554: oled_colour = 16'b00001_001001_00110; 
		2555: oled_colour = 16'b00010_001011_00111; 
		2556: oled_colour = 16'b00110_010000_01001; 
		2557: oled_colour = 16'b00001_001010_00110; 
		2558: oled_colour = 16'b00011_001100_00111; 
		2559: oled_colour = 16'b00100_001101_01000; 
		2560: oled_colour = 16'b00010_001011_00111; 
		2561: oled_colour = 16'b00011_001101_01000; 
		2562: oled_colour = 16'b00101_010100_01101; 
		2563: oled_colour = 16'b00101_010110_10000; 
		2564: oled_colour = 16'b00100_010001_01111; 
		2565: oled_colour = 16'b00011_001110_01110; 
		2566: oled_colour = 16'b00010_001100_01101; 
		2567: oled_colour = 16'b00010_001100_01101; 
		2568: oled_colour = 16'b00010_001100_01101; 
		2569: oled_colour = 16'b00010_001100_01101; 
		2570: oled_colour = 16'b00010_001100_01101; 
		2571: oled_colour = 16'b00010_001100_01101; 
		2572: oled_colour = 16'b00010_001100_01101; 
		2573: oled_colour = 16'b00010_001100_01101; 
		2574: oled_colour = 16'b00010_001100_01101; 
		2575: oled_colour = 16'b00010_001100_01101; 
		2576: oled_colour = 16'b00010_001101_01101; 
		2577: oled_colour = 16'b00110_001111_01011; 
		2578: oled_colour = 16'b00011_000101_00010; 
		2579: oled_colour = 16'b00011_000111_00101; 
		2580: oled_colour = 16'b00010_001001_00111; 
		2581: oled_colour = 16'b00011_001001_00110; 
		2582: oled_colour = 16'b00010_000100_00011; 
		2583: oled_colour = 16'b00100_001010_00111; 
		2584: oled_colour = 16'b01110_011110_01110; 
		2585: oled_colour = 16'b10000_100000_01110; 
		2586: oled_colour = 16'b01111_011111_01110; 
		2587: oled_colour = 16'b10000_100001_01110; 
		2588: oled_colour = 16'b01110_011101_01101; 
		2589: oled_colour = 16'b00110_001111_01000; 
		2590: oled_colour = 16'b01111_011111_01110; 
		2591: oled_colour = 16'b01101_011011_01101; 
		2592: oled_colour = 16'b01001_010010_01000; 
		2593: oled_colour = 16'b00110_001100_00110; 
		2594: oled_colour = 16'b00010_000100_00010; 
		2595: oled_colour = 16'b00010_000101_00100; 
		2596: oled_colour = 16'b00100_001011_01000; 
		2597: oled_colour = 16'b01100_011011_01101; 
		2598: oled_colour = 16'b10110_101100_10001; 
		2599: oled_colour = 16'b11100_110110_10100; 
		2600: oled_colour = 16'b11100_110111_10100; 
		2601: oled_colour = 16'b11000_101110_10010; 
		2602: oled_colour = 16'b01000_010011_01010; 
		2603: oled_colour = 16'b00100_001110_01100; 
		2604: oled_colour = 16'b00011_001110_01101; 
		2605: oled_colour = 16'b00011_001111_01101; 
		2606: oled_colour = 16'b00100_001111_01101; 
		2607: oled_colour = 16'b00100_010000_01101; 
		2608: oled_colour = 16'b00100_010000_01101; 
		2609: oled_colour = 16'b00100_010000_01101; 
		2610: oled_colour = 16'b00100_010000_01101; 
		2611: oled_colour = 16'b00100_010000_01101; 
		2612: oled_colour = 16'b00100_010000_01101; 
		2613: oled_colour = 16'b00100_010000_01101; 
		2614: oled_colour = 16'b00100_010000_01101; 
		2615: oled_colour = 16'b00100_010000_01101; 
		2616: oled_colour = 16'b00100_010000_01101; 
		2617: oled_colour = 16'b00100_010000_01101; 
		2618: oled_colour = 16'b00100_010000_01101; 
		2619: oled_colour = 16'b00100_001111_01101; 
		2620: oled_colour = 16'b00100_001111_01101; 
		2621: oled_colour = 16'b00100_001111_01101; 
		2622: oled_colour = 16'b00100_001111_01101; 
		2623: oled_colour = 16'b00100_010000_01101; 
		2624: oled_colour = 16'b00100_010000_01101; 
		2625: oled_colour = 16'b00100_001111_01101; 
		2626: oled_colour = 16'b00100_010000_01101; 
		2627: oled_colour = 16'b00100_001111_01101; 
		2628: oled_colour = 16'b00100_010000_01101; 
		2629: oled_colour = 16'b00100_010000_01101; 
		2630: oled_colour = 16'b00100_001111_01101; 
		2631: oled_colour = 16'b00100_010000_01101; 
		2632: oled_colour = 16'b00100_001111_01101; 
		2633: oled_colour = 16'b00100_001111_01101; 
		2634: oled_colour = 16'b00100_010000_01101; 
		2635: oled_colour = 16'b00100_010000_01101; 
		2636: oled_colour = 16'b00100_001111_01101; 
		2637: oled_colour = 16'b00100_010001_01110; 
		2638: oled_colour = 16'b01000_011011_10010; 
		2639: oled_colour = 16'b00111_011001_10001; 
		2640: oled_colour = 16'b00111_011000_10000; 
		2641: oled_colour = 16'b00100_001111_01010; 
		2642: oled_colour = 16'b00011_001101_01001; 
		2643: oled_colour = 16'b00010_001010_00111; 
		2644: oled_colour = 16'b00010_001010_00111; 
		2645: oled_colour = 16'b00010_001011_00111; 
		2646: oled_colour = 16'b00010_001010_00110; 
		2647: oled_colour = 16'b00010_001011_00111; 
		2648: oled_colour = 16'b00010_001001_00110; 
		2649: oled_colour = 16'b00001_001000_00101; 
		2650: oled_colour = 16'b00001_001001_00110; 
		2651: oled_colour = 16'b00011_001110_01000; 
		2652: oled_colour = 16'b00011_001101_01000; 
		2653: oled_colour = 16'b00110_010010_01011; 
		2654: oled_colour = 16'b00101_010000_01010; 
		2655: oled_colour = 16'b00011_001100_00111; 
		2656: oled_colour = 16'b00011_001100_00111; 
		2657: oled_colour = 16'b00001_001000_00100; 
		2658: oled_colour = 16'b00001_001010_00110; 
		2659: oled_colour = 16'b00011_001111_01001; 
		2660: oled_colour = 16'b00101_010011_01100; 
		2661: oled_colour = 16'b00110_010110_01111; 
		2662: oled_colour = 16'b01000_011100_10011; 
		2663: oled_colour = 16'b00111_010110_10001; 
		2664: oled_colour = 16'b00100_001111_01101; 
		2665: oled_colour = 16'b00100_010000_01101; 
		2666: oled_colour = 16'b00100_010000_01101; 
		2667: oled_colour = 16'b00100_001111_01101; 
		2668: oled_colour = 16'b00100_010000_01101; 
		2669: oled_colour = 16'b00100_010000_01101; 
		2670: oled_colour = 16'b00100_010000_01101; 
		2671: oled_colour = 16'b00011_001111_01100; 
		2672: oled_colour = 16'b00110_010010_01110; 
		2673: oled_colour = 16'b00110_001100_00111; 
		2674: oled_colour = 16'b00010_000100_00010; 
		2675: oled_colour = 16'b00011_001000_00110; 
		2676: oled_colour = 16'b00010_001001_00111; 
		2677: oled_colour = 16'b00011_000111_00101; 
		2678: oled_colour = 16'b00010_000100_00010; 
		2679: oled_colour = 16'b00010_000111_00101; 
		2680: oled_colour = 16'b01011_011000_01100; 
		2681: oled_colour = 16'b10001_100010_01111; 
		2682: oled_colour = 16'b10000_100001_01110; 
		2683: oled_colour = 16'b10000_100001_01110; 
		2684: oled_colour = 16'b10001_100010_01111; 
		2685: oled_colour = 16'b01001_010101_01010; 
		2686: oled_colour = 16'b01001_010011_01011; 
		2687: oled_colour = 16'b01110_011101_01101; 
		2688: oled_colour = 16'b01000_010010_01001; 
		2689: oled_colour = 16'b00111_010000_01001; 
		2690: oled_colour = 16'b00101_001011_00110; 
		2691: oled_colour = 16'b00010_000101_00011; 
		2692: oled_colour = 16'b00010_000100_00010; 
		2693: oled_colour = 16'b00010_000110_00101; 
		2694: oled_colour = 16'b00110_001110_01000; 
		2695: oled_colour = 16'b01100_011001_01101; 
		2696: oled_colour = 16'b10110_101011_10001; 
		2697: oled_colour = 16'b10111_101101_10001; 
		2698: oled_colour = 16'b01011_011000_01011; 
		2699: oled_colour = 16'b10100_101001_10001; 
		2700: oled_colour = 16'b01100_011100_01110; 
		2701: oled_colour = 16'b00111_010011_01101; 
		2702: oled_colour = 16'b00101_010001_01100; 
		2703: oled_colour = 16'b00100_010000_01101; 
		2704: oled_colour = 16'b00100_010001_01101; 
		2705: oled_colour = 16'b00101_010001_01101; 
		2706: oled_colour = 16'b00100_010001_01101; 
		2707: oled_colour = 16'b00100_010001_01101; 
		2708: oled_colour = 16'b00100_010001_01101; 
		2709: oled_colour = 16'b00100_010001_01101; 
		2710: oled_colour = 16'b00100_010001_01101; 
		2711: oled_colour = 16'b00100_010001_01101; 
		2712: oled_colour = 16'b00100_010001_01101; 
		2713: oled_colour = 16'b00100_010001_01101; 
		2714: oled_colour = 16'b00100_010000_01101; 
		2715: oled_colour = 16'b00100_010000_01101; 
		2716: oled_colour = 16'b00100_010000_01101; 
		2717: oled_colour = 16'b00100_010000_01101; 
		2718: oled_colour = 16'b00100_010000_01101; 
		2719: oled_colour = 16'b00100_010000_01101; 
		2720: oled_colour = 16'b00100_010001_01101; 
		2721: oled_colour = 16'b00100_010001_01101; 
		2722: oled_colour = 16'b00100_010000_01101; 
		2723: oled_colour = 16'b00100_010000_01101; 
		2724: oled_colour = 16'b00100_010000_01101; 
		2725: oled_colour = 16'b00100_010000_01101; 
		2726: oled_colour = 16'b00100_010001_01101; 
		2727: oled_colour = 16'b00100_010001_01101; 
		2728: oled_colour = 16'b00100_010000_01101; 
		2729: oled_colour = 16'b00100_010000_01101; 
		2730: oled_colour = 16'b00100_010000_01101; 
		2731: oled_colour = 16'b00100_010001_01101; 
		2732: oled_colour = 16'b00100_010000_01100; 
		2733: oled_colour = 16'b00110_010100_01111; 
		2734: oled_colour = 16'b00110_010100_01101; 
		2735: oled_colour = 16'b00011_001110_01001; 
		2736: oled_colour = 16'b00011_001101_01000; 
		2737: oled_colour = 16'b00001_000100_00011; 
		2738: oled_colour = 16'b00001_000100_00010; 
		2739: oled_colour = 16'b00001_000110_00100; 
		2740: oled_colour = 16'b00001_000111_00101; 
		2741: oled_colour = 16'b00001_000111_00101; 
		2742: oled_colour = 16'b00010_001001_00101; 
		2743: oled_colour = 16'b00011_001010_00110; 
		2744: oled_colour = 16'b00010_001010_00110; 
		2745: oled_colour = 16'b00010_001011_00111; 
		2746: oled_colour = 16'b00011_001100_00111; 
		2747: oled_colour = 16'b00100_001110_01001; 
		2748: oled_colour = 16'b00100_001111_01001; 
		2749: oled_colour = 16'b00100_001100_01000; 
		2750: oled_colour = 16'b00101_001111_01010; 
		2751: oled_colour = 16'b00100_001111_01001; 
		2752: oled_colour = 16'b00011_001101_00111; 
		2753: oled_colour = 16'b00101_001101_00111; 
		2754: oled_colour = 16'b00011_001001_00110; 
		2755: oled_colour = 16'b00010_001000_00101; 
		2756: oled_colour = 16'b00001_000110_00100; 
		2757: oled_colour = 16'b00010_001100_01000; 
		2758: oled_colour = 16'b00111_011000_10000; 
		2759: oled_colour = 16'b00101_010011_01110; 
		2760: oled_colour = 16'b00100_010000_01101; 
		2761: oled_colour = 16'b00100_010001_01101; 
		2762: oled_colour = 16'b00100_010001_01101; 
		2763: oled_colour = 16'b00100_010000_01101; 
		2764: oled_colour = 16'b00100_010000_01101; 
		2765: oled_colour = 16'b00100_010000_01101; 
		2766: oled_colour = 16'b00100_010000_01100; 
		2767: oled_colour = 16'b00100_010001_01101; 
		2768: oled_colour = 16'b01000_010100_01110; 
		2769: oled_colour = 16'b00100_000110_00011; 
		2770: oled_colour = 16'b00010_000110_00100; 
		2771: oled_colour = 16'b00010_001001_00111; 
		2772: oled_colour = 16'b00011_001001_00111; 
		2773: oled_colour = 16'b00011_000110_00011; 
		2774: oled_colour = 16'b00011_000101_00010; 
		2775: oled_colour = 16'b00010_000101_00100; 
		2776: oled_colour = 16'b01010_010110_01100; 
		2777: oled_colour = 16'b01110_011101_01110; 
		2778: oled_colour = 16'b01101_011010_01100; 
		2779: oled_colour = 16'b01101_011011_01101; 
		2780: oled_colour = 16'b01100_011000_01100; 
		2781: oled_colour = 16'b01010_010111_01010; 
		2782: oled_colour = 16'b00111_010001_01001; 
		2783: oled_colour = 16'b10010_100101_10000; 
		2784: oled_colour = 16'b00111_010010_01011; 
		2785: oled_colour = 16'b00011_001001_00110; 
		2786: oled_colour = 16'b00100_001011_00111; 
		2787: oled_colour = 16'b00100_001010_00110; 
		2788: oled_colour = 16'b00010_000101_00011; 
		2789: oled_colour = 16'b00010_000100_00010; 
		2790: oled_colour = 16'b00010_000100_00010; 
		2791: oled_colour = 16'b00010_000110_00101; 
		2792: oled_colour = 16'b00110_001111_01001; 
		2793: oled_colour = 16'b00110_001110_01000; 
		2794: oled_colour = 16'b01010_010110_01100; 
		2795: oled_colour = 16'b11001_110001_10011; 
		2796: oled_colour = 16'b11100_110110_10011; 
		2797: oled_colour = 16'b10110_101100_10001; 
		2798: oled_colour = 16'b01111_100001_01110; 
		2799: oled_colour = 16'b01011_011010_01110; 
		2800: oled_colour = 16'b00110_010011_01101; 
		2801: oled_colour = 16'b00101_010010_01110; 
		2802: oled_colour = 16'b00110_010011_01110; 
		2803: oled_colour = 16'b00110_010011_01110; 
		2804: oled_colour = 16'b00101_010011_01110; 
		2805: oled_colour = 16'b00110_010011_01110; 
		2806: oled_colour = 16'b00110_010011_01110; 
		2807: oled_colour = 16'b00101_010011_01110; 
		2808: oled_colour = 16'b00101_010011_01110; 
		2809: oled_colour = 16'b00110_010011_01110; 
		2810: oled_colour = 16'b00101_010011_01110; 
		2811: oled_colour = 16'b00101_010011_01110; 
		2812: oled_colour = 16'b00101_010011_01110; 
		2813: oled_colour = 16'b00101_010011_01110; 
		2814: oled_colour = 16'b00101_010011_01110; 
		2815: oled_colour = 16'b00110_010011_01110; 
		2816: oled_colour = 16'b00101_010011_01110; 
		2817: oled_colour = 16'b00110_010011_01110; 
		2818: oled_colour = 16'b00110_010011_01110; 
		2819: oled_colour = 16'b00101_010011_01110; 
		2820: oled_colour = 16'b00101_010011_01110; 
		2821: oled_colour = 16'b00101_010011_01110; 
		2822: oled_colour = 16'b00101_010011_01110; 
		2823: oled_colour = 16'b00101_010011_01110; 
		2824: oled_colour = 16'b00101_010011_01110; 
		2825: oled_colour = 16'b00101_010011_01110; 
		2826: oled_colour = 16'b00101_010011_01110; 
		2827: oled_colour = 16'b00110_010011_01110; 
		2828: oled_colour = 16'b00101_010010_01110; 
		2829: oled_colour = 16'b00111_010111_10001; 
		2830: oled_colour = 16'b00101_010011_01100; 
		2831: oled_colour = 16'b00001_001001_00101; 
		2832: oled_colour = 16'b00001_000110_00100; 
		2833: oled_colour = 16'b00001_000100_00011; 
		2834: oled_colour = 16'b00001_000101_00100; 
		2835: oled_colour = 16'b00111_010010_01010; 
		2836: oled_colour = 16'b00011_001011_00111; 
		2837: oled_colour = 16'b00001_000011_00010; 
		2838: oled_colour = 16'b00011_001010_00110; 
		2839: oled_colour = 16'b00100_001101_01000; 
		2840: oled_colour = 16'b00010_001011_00111; 
		2841: oled_colour = 16'b00010_001011_00111; 
		2842: oled_colour = 16'b00100_010000_01010; 
		2843: oled_colour = 16'b00111_010011_01101; 
		2844: oled_colour = 16'b00011_001101_01001; 
		2845: oled_colour = 16'b00001_001000_00110; 
		2846: oled_colour = 16'b00010_001011_01000; 
		2847: oled_colour = 16'b00111_010011_01100; 
		2848: oled_colour = 16'b00100_010000_01010; 
		2849: oled_colour = 16'b00011_001100_00111; 
		2850: oled_colour = 16'b00100_001101_01000; 
		2851: oled_colour = 16'b00100_001101_01000; 
		2852: oled_colour = 16'b00100_001110_01001; 
		2853: oled_colour = 16'b00110_010110_01110; 
		2854: oled_colour = 16'b00110_010101_01111; 
		2855: oled_colour = 16'b00101_010010_01101; 
		2856: oled_colour = 16'b00110_010011_01110; 
		2857: oled_colour = 16'b00101_010010_01110; 
		2858: oled_colour = 16'b00101_010011_01110; 
		2859: oled_colour = 16'b00101_010011_01110; 
		2860: oled_colour = 16'b00101_010011_01110; 
		2861: oled_colour = 16'b00101_010010_01110; 
		2862: oled_colour = 16'b00101_010010_01110; 
		2863: oled_colour = 16'b00110_010100_01111; 
		2864: oled_colour = 16'b00111_001111_01010; 
		2865: oled_colour = 16'b00010_000100_00010; 
		2866: oled_colour = 16'b00011_001000_00110; 
		2867: oled_colour = 16'b00010_001001_00111; 
		2868: oled_colour = 16'b00011_001000_00101; 
		2869: oled_colour = 16'b00010_000100_00010; 
		2870: oled_colour = 16'b00011_000101_00011; 
		2871: oled_colour = 16'b00010_000101_00011; 
		2872: oled_colour = 16'b00100_001100_01000; 
		2873: oled_colour = 16'b10000_100001_01110; 
		2874: oled_colour = 16'b10001_100001_01110; 
		2875: oled_colour = 16'b10001_100011_01111; 
		2876: oled_colour = 16'b10001_100010_01110; 
		2877: oled_colour = 16'b01111_100000_01110; 
		2878: oled_colour = 16'b00101_001110_01000; 
		2879: oled_colour = 16'b10000_100000_01110; 
		2880: oled_colour = 16'b00011_001000_00101; 
		2881: oled_colour = 16'b00101_001101_01000; 
		2882: oled_colour = 16'b01011_011000_01100; 
		2883: oled_colour = 16'b00101_001101_01000; 
		2884: oled_colour = 16'b00011_001001_00111; 
		2885: oled_colour = 16'b00011_000110_00101; 
		2886: oled_colour = 16'b00011_000101_00011; 
		2887: oled_colour = 16'b00011_000101_00011; 
		2888: oled_colour = 16'b00010_000100_00011; 
		2889: oled_colour = 16'b00010_000100_00011; 
		2890: oled_colour = 16'b00100_001001_00111; 
		2891: oled_colour = 16'b01000_010011_01011; 
		2892: oled_colour = 16'b10010_100100_10000; 
		2893: oled_colour = 16'b11001_110010_10010; 
		2894: oled_colour = 16'b11101_111000_10100; 
		2895: oled_colour = 16'b10101_101011_10000; 
		2896: oled_colour = 16'b00111_010001_01010; 
		2897: oled_colour = 16'b01000_010110_01111; 
		2898: oled_colour = 16'b00111_010100_10000; 
		2899: oled_colour = 16'b00111_010101_10000; 
		2900: oled_colour = 16'b00111_010101_10000; 
		2901: oled_colour = 16'b00111_010101_10000; 
		2902: oled_colour = 16'b00111_010101_10000; 
		2903: oled_colour = 16'b00111_010101_10000; 
		2904: oled_colour = 16'b00111_010101_01111; 
		2905: oled_colour = 16'b00111_010101_10000; 
		2906: oled_colour = 16'b00111_010101_10000; 
		2907: oled_colour = 16'b00111_010101_10000; 
		2908: oled_colour = 16'b00111_010101_10000; 
		2909: oled_colour = 16'b00111_010101_10000; 
		2910: oled_colour = 16'b00111_010101_10000; 
		2911: oled_colour = 16'b00111_010101_10000; 
		2912: oled_colour = 16'b00111_010101_10000; 
		2913: oled_colour = 16'b00111_010101_10000; 
		2914: oled_colour = 16'b00111_010101_10000; 
		2915: oled_colour = 16'b00111_010101_10000; 
		2916: oled_colour = 16'b00111_010101_10000; 
		2917: oled_colour = 16'b00111_010101_01111; 
		2918: oled_colour = 16'b00111_010101_01111; 
		2919: oled_colour = 16'b00111_010101_01111; 
		2920: oled_colour = 16'b00111_010101_10000; 
		2921: oled_colour = 16'b00111_010101_10000; 
		2922: oled_colour = 16'b00111_010101_10000; 
		2923: oled_colour = 16'b00111_010101_10000; 
		2924: oled_colour = 16'b00111_010101_01111; 
		2925: oled_colour = 16'b01000_011001_10001; 
		2926: oled_colour = 16'b00100_010000_01010; 
		2927: oled_colour = 16'b00001_000111_00100; 
		2928: oled_colour = 16'b00001_000100_00011; 
		2929: oled_colour = 16'b00001_000100_00011; 
		2930: oled_colour = 16'b00010_001010_00110; 
		2931: oled_colour = 16'b00101_010001_01010; 
		2932: oled_colour = 16'b00010_001001_00110; 
		2933: oled_colour = 16'b00100_001101_01000; 
		2934: oled_colour = 16'b00110_010000_01010; 
		2935: oled_colour = 16'b00101_001111_01001; 
		2936: oled_colour = 16'b00011_001100_01000; 
		2937: oled_colour = 16'b00010_001011_00111; 
		2938: oled_colour = 16'b00011_001101_01001; 
		2939: oled_colour = 16'b00011_001110_01001; 
		2940: oled_colour = 16'b00011_001101_01001; 
		2941: oled_colour = 16'b00011_001101_01001; 
		2942: oled_colour = 16'b00011_001100_01000; 
		2943: oled_colour = 16'b00011_001101_01000; 
		2944: oled_colour = 16'b00011_001100_01000; 
		2945: oled_colour = 16'b00011_001100_01000; 
		2946: oled_colour = 16'b00011_001100_01000; 
		2947: oled_colour = 16'b00100_001110_01001; 
		2948: oled_colour = 16'b00110_010010_01011; 
		2949: oled_colour = 16'b01000_010100_01100; 
		2950: oled_colour = 16'b00111_010011_01100; 
		2951: oled_colour = 16'b00111_010101_10000; 
		2952: oled_colour = 16'b00111_010101_10000; 
		2953: oled_colour = 16'b00111_010101_10000; 
		2954: oled_colour = 16'b00111_010101_10000; 
		2955: oled_colour = 16'b00111_010101_10000; 
		2956: oled_colour = 16'b00111_010101_10000; 
		2957: oled_colour = 16'b00111_010101_10000; 
		2958: oled_colour = 16'b00111_010101_01111; 
		2959: oled_colour = 16'b01010_011000_10000; 
		2960: oled_colour = 16'b00100_000111_00100; 
		2961: oled_colour = 16'b00010_000100_00011; 
		2962: oled_colour = 16'b00010_001001_00111; 
		2963: oled_colour = 16'b00010_001001_00111; 
		2964: oled_colour = 16'b00011_000110_00100; 
		2965: oled_colour = 16'b00011_000100_00010; 
		2966: oled_colour = 16'b00011_000101_00011; 
		2967: oled_colour = 16'b00010_000100_00010; 
		2968: oled_colour = 16'b00011_001000_00110; 
		2969: oled_colour = 16'b01100_011001_01101; 
		2970: oled_colour = 16'b01110_011101_01101; 
		2971: oled_colour = 16'b10000_011111_01110; 
		2972: oled_colour = 16'b10000_011111_01110; 
		2973: oled_colour = 16'b10000_100010_01110; 
		2974: oled_colour = 16'b01100_011011_01100; 
		2975: oled_colour = 16'b01010_010100_01010; 
		2976: oled_colour = 16'b00101_001101_01000; 
		2977: oled_colour = 16'b00101_001101_01000; 
		2978: oled_colour = 16'b00101_001101_01001; 
		2979: oled_colour = 16'b00011_000111_00110; 
		2980: oled_colour = 16'b00100_001001_00111; 
		2981: oled_colour = 16'b00010_000101_00100; 
		2982: oled_colour = 16'b00011_000110_00101; 
		2983: oled_colour = 16'b00011_000110_00100; 
		2984: oled_colour = 16'b00011_000101_00011; 
		2985: oled_colour = 16'b00011_000101_00011; 
		2986: oled_colour = 16'b00010_000100_00010; 
		2987: oled_colour = 16'b00010_000101_00100; 
		2988: oled_colour = 16'b00100_001010_01000; 
		2989: oled_colour = 16'b01001_010101_01011; 
		2990: oled_colour = 16'b10110_101011_10010; 
		2991: oled_colour = 16'b10000_100001_01110; 
		2992: oled_colour = 16'b10001_100100_01111; 
		2993: oled_colour = 16'b11000_110000_10010; 
		2994: oled_colour = 16'b01111_100001_10000; 
		2995: oled_colour = 16'b01011_011010_10000; 
		2996: oled_colour = 16'b01010_011000_10001; 
		2997: oled_colour = 16'b01010_011000_10010; 
		2998: oled_colour = 16'b01010_011001_10010; 
		2999: oled_colour = 16'b01010_011001_10010; 
		3000: oled_colour = 16'b01010_011001_10001; 
		3001: oled_colour = 16'b01010_011000_10010; 
		3002: oled_colour = 16'b01010_011000_10010; 
		3003: oled_colour = 16'b01010_011000_10010; 
		3004: oled_colour = 16'b01010_011001_10010; 
		3005: oled_colour = 16'b01010_011001_10010; 
		3006: oled_colour = 16'b01010_011001_10010; 
		3007: oled_colour = 16'b01010_011001_10010; 
		3008: oled_colour = 16'b01010_011001_10010; 
		3009: oled_colour = 16'b01010_011001_10001; 
		3010: oled_colour = 16'b01010_011001_10010; 
		3011: oled_colour = 16'b01010_011001_10010; 
		3012: oled_colour = 16'b01010_011001_10010; 
		3013: oled_colour = 16'b01010_011001_10010; 
		3014: oled_colour = 16'b01010_011001_10010; 
		3015: oled_colour = 16'b01010_011000_10010; 
		3016: oled_colour = 16'b01010_011001_10010; 
		3017: oled_colour = 16'b01010_011000_10010; 
		3018: oled_colour = 16'b01010_011001_10010; 
		3019: oled_colour = 16'b01010_011000_10010; 
		3020: oled_colour = 16'b01010_011000_10010; 
		3021: oled_colour = 16'b01001_011010_10001; 
		3022: oled_colour = 16'b00010_001011_00111; 
		3023: oled_colour = 16'b00001_000110_00100; 
		3024: oled_colour = 16'b00001_000101_00011; 
		3025: oled_colour = 16'b00001_000100_00011; 
		3026: oled_colour = 16'b00010_001011_00111; 
		3027: oled_colour = 16'b00001_001011_00111; 
		3028: oled_colour = 16'b00001_000100_00011; 
		3029: oled_colour = 16'b00001_000110_00100; 
		3030: oled_colour = 16'b00010_000111_00100; 
		3031: oled_colour = 16'b00011_001001_00101; 
		3032: oled_colour = 16'b00011_001010_00110; 
		3033: oled_colour = 16'b00011_001010_00110; 
		3034: oled_colour = 16'b00010_001001_00101; 
		3035: oled_colour = 16'b00011_001010_00110; 
		3036: oled_colour = 16'b00010_001001_00101; 
		3037: oled_colour = 16'b00010_001001_00101; 
		3038: oled_colour = 16'b00011_001001_00101; 
		3039: oled_colour = 16'b00010_001001_00101; 
		3040: oled_colour = 16'b00010_001000_00101; 
		3041: oled_colour = 16'b00011_001001_00101; 
		3042: oled_colour = 16'b00011_001010_00110; 
		3043: oled_colour = 16'b00011_001010_00110; 
		3044: oled_colour = 16'b00010_001000_00101; 
		3045: oled_colour = 16'b00010_001000_00101; 
		3046: oled_colour = 16'b00111_010011_01101; 
		3047: oled_colour = 16'b01010_011001_10010; 
		3048: oled_colour = 16'b01010_011001_10001; 
		3049: oled_colour = 16'b01010_011001_10010; 
		3050: oled_colour = 16'b01010_011001_10010; 
		3051: oled_colour = 16'b01010_011000_10010; 
		3052: oled_colour = 16'b01010_011000_10010; 
		3053: oled_colour = 16'b01010_011000_10001; 
		3054: oled_colour = 16'b01011_011011_10011; 
		3055: oled_colour = 16'b01000_010000_01010; 
		3056: oled_colour = 16'b00010_000011_00001; 
		3057: oled_colour = 16'b00011_000101_00011; 
		3058: oled_colour = 16'b00010_001000_00111; 
		3059: oled_colour = 16'b00011_001001_00110; 
		3060: oled_colour = 16'b00011_000101_00011; 
		3061: oled_colour = 16'b00011_000101_00010; 
		3062: oled_colour = 16'b00011_000101_00011; 
		3063: oled_colour = 16'b00011_000101_00010; 
		3064: oled_colour = 16'b00010_000101_00100; 
		3065: oled_colour = 16'b01001_010100_01011; 
		3066: oled_colour = 16'b10010_100100_10000; 
		3067: oled_colour = 16'b01111_011110_01101; 
		3068: oled_colour = 16'b01111_011101_01101; 
		3069: oled_colour = 16'b01110_011100_01101; 
		3070: oled_colour = 16'b01010_010110_01011; 
		3071: oled_colour = 16'b00110_001110_01000; 
		3072: oled_colour = 16'b00101_001100_01000; 
		3073: oled_colour = 16'b00101_001100_01000; 
		3074: oled_colour = 16'b00101_001101_01000; 
		3075: oled_colour = 16'b00110_001101_01000; 
		3076: oled_colour = 16'b00100_001001_00111; 
		3077: oled_colour = 16'b00011_000101_00011; 
		3078: oled_colour = 16'b00011_000101_00011; 
		3079: oled_colour = 16'b00011_000101_00100; 
		3080: oled_colour = 16'b00011_000110_00101; 
		3081: oled_colour = 16'b00011_000111_00101; 
		3082: oled_colour = 16'b00011_000110_00011; 
		3083: oled_colour = 16'b00011_000101_00010; 
		3084: oled_colour = 16'b00010_000100_00010; 
		3085: oled_colour = 16'b00010_000101_00100; 
		3086: oled_colour = 16'b00100_001010_00111; 
		3087: oled_colour = 16'b00100_001010_00110; 
		3088: oled_colour = 16'b01010_010111_01011; 
		3089: oled_colour = 16'b10110_101100_10001; 
		3090: oled_colour = 16'b11100_110111_10011; 
		3091: oled_colour = 16'b11010_110010_10010; 
		3092: oled_colour = 16'b10100_101001_10000; 
		3093: oled_colour = 16'b01110_100000_01111; 
		3094: oled_colour = 16'b01100_011100_10000; 
		3095: oled_colour = 16'b01011_011010_10001; 
		3096: oled_colour = 16'b01100_011011_10010; 
		3097: oled_colour = 16'b01100_011100_10010; 
		3098: oled_colour = 16'b01011_011011_10010; 
		3099: oled_colour = 16'b01100_011011_10010; 
		3100: oled_colour = 16'b01100_011011_10010; 
		3101: oled_colour = 16'b01100_011011_10010; 
		3102: oled_colour = 16'b01100_011011_10010; 
		3103: oled_colour = 16'b01100_011011_10010; 
		3104: oled_colour = 16'b01100_011011_10010; 
		3105: oled_colour = 16'b01100_011100_10010; 
		3106: oled_colour = 16'b01011_011100_10010; 
		3107: oled_colour = 16'b01100_011011_10010; 
		3108: oled_colour = 16'b01100_011011_10010; 
		3109: oled_colour = 16'b01011_011011_10010; 
		3110: oled_colour = 16'b01100_011011_10010; 
		3111: oled_colour = 16'b01100_011011_10010; 
		3112: oled_colour = 16'b01100_011011_10010; 
		3113: oled_colour = 16'b01100_011011_10010; 
		3114: oled_colour = 16'b01100_011011_10010; 
		3115: oled_colour = 16'b01100_011011_10010; 
		3116: oled_colour = 16'b01100_011100_10010; 
		3117: oled_colour = 16'b01010_011100_10001; 
		3118: oled_colour = 16'b00001_001000_00101; 
		3119: oled_colour = 16'b00010_001001_00101; 
		3120: oled_colour = 16'b00001_001000_00101; 
		3121: oled_colour = 16'b00001_000111_00100; 
		3122: oled_colour = 16'b00010_001010_00110; 
		3123: oled_colour = 16'b00011_001101_01000; 
		3124: oled_colour = 16'b00010_000111_00100; 
		3125: oled_colour = 16'b00001_000101_00011; 
		3126: oled_colour = 16'b00010_001010_00110; 
		3127: oled_colour = 16'b00010_001011_00111; 
		3128: oled_colour = 16'b00010_001001_00101; 
		3129: oled_colour = 16'b00010_001100_00111; 
		3130: oled_colour = 16'b00010_001100_00111; 
		3131: oled_colour = 16'b00010_001001_00110; 
		3132: oled_colour = 16'b00001_001000_00101; 
		3133: oled_colour = 16'b00001_000100_00011; 
		3134: oled_colour = 16'b00001_000111_00100; 
		3135: oled_colour = 16'b00010_001001_00110; 
		3136: oled_colour = 16'b00001_001001_00110; 
		3137: oled_colour = 16'b00010_001000_00101; 
		3138: oled_colour = 16'b00001_000111_00100; 
		3139: oled_colour = 16'b00001_000111_00100; 
		3140: oled_colour = 16'b00011_001010_00111; 
		3141: oled_colour = 16'b00100_010001_01010; 
		3142: oled_colour = 16'b01011_100000_10100; 
		3143: oled_colour = 16'b01100_011100_10010; 
		3144: oled_colour = 16'b01100_011011_10010; 
		3145: oled_colour = 16'b01100_011011_10010; 
		3146: oled_colour = 16'b01011_011011_10010; 
		3147: oled_colour = 16'b01100_011011_10010; 
		3148: oled_colour = 16'b01100_011011_10010; 
		3149: oled_colour = 16'b01100_011101_10011; 
		3150: oled_colour = 16'b01100_011010_10000; 
		3151: oled_colour = 16'b00011_000110_00011; 
		3152: oled_colour = 16'b00011_000101_00011; 
		3153: oled_colour = 16'b00011_000110_00100; 
		3154: oled_colour = 16'b00011_001001_00111; 
		3155: oled_colour = 16'b00011_001000_00101; 
		3156: oled_colour = 16'b00011_000101_00010; 
		3157: oled_colour = 16'b00011_000101_00011; 
		3158: oled_colour = 16'b00011_000101_00011; 
		3159: oled_colour = 16'b00011_000101_00011; 
		3160: oled_colour = 16'b00010_000101_00011; 
		3161: oled_colour = 16'b00101_001100_01000; 
		3162: oled_colour = 16'b01010_010110_01011; 
		3163: oled_colour = 16'b01101_011011_01101; 
		3164: oled_colour = 16'b01110_011101_01101; 
		3165: oled_colour = 16'b10000_100000_01110; 
		3166: oled_colour = 16'b10010_100100_01111; 
		3167: oled_colour = 16'b01000_010011_01001; 
		3168: oled_colour = 16'b01001_010101_01100; 
		3169: oled_colour = 16'b00100_001011_01000; 
		3170: oled_colour = 16'b00110_001110_01001; 
		3171: oled_colour = 16'b00111_010000_01010; 
		3172: oled_colour = 16'b00100_001011_01000; 
		3173: oled_colour = 16'b00011_000110_00100; 
		3174: oled_colour = 16'b00010_000100_00010; 
		3175: oled_colour = 16'b00011_000101_00011; 
		3176: oled_colour = 16'b00010_000101_00011; 
		3177: oled_colour = 16'b00010_000101_00100; 
		3178: oled_colour = 16'b00011_000110_00100; 
		3179: oled_colour = 16'b00011_000110_00101; 
		3180: oled_colour = 16'b00011_000110_00100; 
		3181: oled_colour = 16'b00011_000101_00010; 
		3182: oled_colour = 16'b00010_000100_00010; 
		3183: oled_colour = 16'b00010_000100_00010; 
		3184: oled_colour = 16'b00010_000100_00011; 
		3185: oled_colour = 16'b00100_001010_00110; 
		3186: oled_colour = 16'b01101_011010_01101; 
		3187: oled_colour = 16'b10111_101110_10010; 
		3188: oled_colour = 16'b11100_110111_10100; 
		3189: oled_colour = 16'b11100_110110_10011; 
		3190: oled_colour = 16'b10110_101011_10000; 
		3191: oled_colour = 16'b01001_010100_01011; 
		3192: oled_colour = 16'b01101_011100_10000; 
		3193: oled_colour = 16'b01111_011111_10010; 
		3194: oled_colour = 16'b10000_100001_10010; 
		3195: oled_colour = 16'b10000_100000_10010; 
		3196: oled_colour = 16'b01111_011111_10010; 
		3197: oled_colour = 16'b01111_011111_10001; 
		3198: oled_colour = 16'b01111_011111_10001; 
		3199: oled_colour = 16'b01111_011111_10001; 
		3200: oled_colour = 16'b01111_011111_10001; 
		3201: oled_colour = 16'b01111_011111_10001; 
		3202: oled_colour = 16'b01111_011111_10001; 
		3203: oled_colour = 16'b01111_011111_10010; 
		3204: oled_colour = 16'b01111_011111_10010; 
		3205: oled_colour = 16'b01111_011111_10001; 
		3206: oled_colour = 16'b01111_011111_10001; 
		3207: oled_colour = 16'b01111_011111_10001; 
		3208: oled_colour = 16'b01111_011111_10001; 
		3209: oled_colour = 16'b01111_011111_10001; 
		3210: oled_colour = 16'b01111_011111_10001; 
		3211: oled_colour = 16'b01111_011111_10001; 
		3212: oled_colour = 16'b10000_100000_10010; 
		3213: oled_colour = 16'b01010_011010_01111; 
		3214: oled_colour = 16'b00001_000001_00010; 
		3215: oled_colour = 16'b00001_000110_00100; 
		3216: oled_colour = 16'b00001_000111_00100; 
		3217: oled_colour = 16'b00001_000101_00011; 
		3218: oled_colour = 16'b00001_000100_00011; 
		3219: oled_colour = 16'b00001_000100_00011; 
		3220: oled_colour = 16'b00001_000011_00010; 
		3221: oled_colour = 16'b00001_000011_00010; 
		3222: oled_colour = 16'b00010_001100_01001; 
		3223: oled_colour = 16'b00010_001101_01001; 
		3224: oled_colour = 16'b00001_000110_00101; 
		3225: oled_colour = 16'b00010_001101_01010; 
		3226: oled_colour = 16'b00011_001110_01010; 
		3227: oled_colour = 16'b00011_001110_01010; 
		3228: oled_colour = 16'b00001_001010_00111; 
		3229: oled_colour = 16'b00001_000011_00010; 
		3230: oled_colour = 16'b00001_001000_00110; 
		3231: oled_colour = 16'b00010_001110_01010; 
		3232: oled_colour = 16'b00010_001110_01010; 
		3233: oled_colour = 16'b00011_001101_01010; 
		3234: oled_colour = 16'b00001_000110_00101; 
		3235: oled_colour = 16'b00001_000111_00101; 
		3236: oled_colour = 16'b00010_001101_01001; 
		3237: oled_colour = 16'b00001_000101_00100; 
		3238: oled_colour = 16'b00101_010101_01101; 
		3239: oled_colour = 16'b01110_100011_10101; 
		3240: oled_colour = 16'b01111_011111_10001; 
		3241: oled_colour = 16'b01111_011111_10001; 
		3242: oled_colour = 16'b01111_011111_10001; 
		3243: oled_colour = 16'b01111_011111_10001; 
		3244: oled_colour = 16'b01111_011111_10001; 
		3245: oled_colour = 16'b01111_100000_10010; 
		3246: oled_colour = 16'b00110_001101_01000; 
		3247: oled_colour = 16'b00001_000001_00001; 
		3248: oled_colour = 16'b00001_000010_00010; 
		3249: oled_colour = 16'b00001_000010_00010; 
		3250: oled_colour = 16'b00001_000110_00101; 
		3251: oled_colour = 16'b00001_000010_00010; 
		3252: oled_colour = 16'b00010_000011_00010; 
		3253: oled_colour = 16'b00010_000100_00010; 
		3254: oled_colour = 16'b00010_000100_00010; 
		3255: oled_colour = 16'b00010_000100_00010; 
		3256: oled_colour = 16'b00010_000100_00010; 
		3257: oled_colour = 16'b00011_001000_00110; 
		3258: oled_colour = 16'b01101_011100_01101; 
		3259: oled_colour = 16'b01111_011110_01110; 
		3260: oled_colour = 16'b01110_011101_01101; 
		3261: oled_colour = 16'b01101_011011_01100; 
		3262: oled_colour = 16'b01100_011001_01100; 
		3263: oled_colour = 16'b01010_010111_01011; 
		3264: oled_colour = 16'b00111_010001_01011; 
		3265: oled_colour = 16'b00011_000111_00101; 
		3266: oled_colour = 16'b00011_001000_00101; 
		3267: oled_colour = 16'b00011_000111_00101; 
		3268: oled_colour = 16'b00101_001100_01001; 
		3269: oled_colour = 16'b00011_000111_00100; 
		3270: oled_colour = 16'b00010_000100_00010; 
		3271: oled_colour = 16'b00011_000101_00011; 
		3272: oled_colour = 16'b00011_000101_00010; 
		3273: oled_colour = 16'b00011_000100_00011; 
		3274: oled_colour = 16'b00011_000100_00011; 
		3275: oled_colour = 16'b00011_000101_00100; 
		3276: oled_colour = 16'b00011_000110_00101; 
		3277: oled_colour = 16'b00011_000111_00101; 
		3278: oled_colour = 16'b00011_000110_00100; 
		3279: oled_colour = 16'b00010_000011_00010; 
		3280: oled_colour = 16'b00010_000010_00010; 
		3281: oled_colour = 16'b00001_000010_00010; 
		3282: oled_colour = 16'b00001_000010_00010; 
		3283: oled_colour = 16'b00100_001010_00110; 
		3284: oled_colour = 16'b01100_011000_01100; 
		3285: oled_colour = 16'b10111_101101_10010; 
		3286: oled_colour = 16'b10101_101001_10000; 
		3287: oled_colour = 16'b01111_011111_01101; 
		3288: oled_colour = 16'b10111_101110_10010; 
		3289: oled_colour = 16'b10001_100010_10000; 
		3290: oled_colour = 16'b10000_100001_10001; 
		3291: oled_colour = 16'b10011_100110_10100; 
		3292: oled_colour = 16'b10101_101010_10101; 
		3293: oled_colour = 16'b10110_101010_10101; 
		3294: oled_colour = 16'b10110_101011_10110; 
		3295: oled_colour = 16'b10110_101011_10110; 
		3296: oled_colour = 16'b10110_101011_10110; 
		3297: oled_colour = 16'b10110_101011_10110; 
		3298: oled_colour = 16'b10110_101011_10110; 
		3299: oled_colour = 16'b10110_101011_10110; 
		3300: oled_colour = 16'b10110_101011_10110; 
		3301: oled_colour = 16'b10110_101011_10110; 
		3302: oled_colour = 16'b10110_101010_10101; 
		3303: oled_colour = 16'b10110_101010_10110; 
		3304: oled_colour = 16'b10110_101010_10110; 
		3305: oled_colour = 16'b10110_101011_10110; 
		3306: oled_colour = 16'b10110_101011_10110; 
		3307: oled_colour = 16'b10110_101010_10110; 
		3308: oled_colour = 16'b10110_101011_10110; 
		3309: oled_colour = 16'b10011_100111_10100; 
		3310: oled_colour = 16'b01110_011101_10000; 
		3311: oled_colour = 16'b01111_011111_10000; 
		3312: oled_colour = 16'b01111_100000_10001; 
		3313: oled_colour = 16'b01111_011111_10000; 
		3314: oled_colour = 16'b01111_011111_10000; 
		3315: oled_colour = 16'b01111_011101_01111; 
		3316: oled_colour = 16'b01111_011101_01111; 
		3317: oled_colour = 16'b01111_011110_01111; 
		3318: oled_colour = 16'b01111_100000_10001; 
		3319: oled_colour = 16'b10000_100001_10010; 
		3320: oled_colour = 16'b01111_011111_10001; 
		3321: oled_colour = 16'b01111_100001_10010; 
		3322: oled_colour = 16'b10000_100001_10010; 
		3323: oled_colour = 16'b10000_100001_10010; 
		3324: oled_colour = 16'b01111_100001_10010; 
		3325: oled_colour = 16'b01111_100000_10001; 
		3326: oled_colour = 16'b01111_100000_10001; 
		3327: oled_colour = 16'b10000_100010_10010; 
		3328: oled_colour = 16'b10000_100010_10010; 
		3329: oled_colour = 16'b10000_100010_10011; 
		3330: oled_colour = 16'b01111_011111_10001; 
		3331: oled_colour = 16'b01111_011111_10001; 
		3332: oled_colour = 16'b10000_100010_10010; 
		3333: oled_colour = 16'b01111_011110_10000; 
		3334: oled_colour = 16'b01111_100001_10010; 
		3335: oled_colour = 16'b10100_101100_11000; 
		3336: oled_colour = 16'b10110_101011_10110; 
		3337: oled_colour = 16'b10110_101011_10110; 
		3338: oled_colour = 16'b10110_101011_10110; 
		3339: oled_colour = 16'b10110_101011_10110; 
		3340: oled_colour = 16'b10110_101011_10110; 
		3341: oled_colour = 16'b10101_101000_10101; 
		3342: oled_colour = 16'b01111_011110_01111; 
		3343: oled_colour = 16'b01111_011110_01111; 
		3344: oled_colour = 16'b01111_011110_01111; 
		3345: oled_colour = 16'b01111_011110_10000; 
		3346: oled_colour = 16'b10000_100000_10001; 
		3347: oled_colour = 16'b10000_100000_10000; 
		3348: oled_colour = 16'b01001_010011_01001; 
		3349: oled_colour = 16'b00101_001010_00111; 
		3350: oled_colour = 16'b00101_001011_00111; 
		3351: oled_colour = 16'b00100_001010_00110; 
		3352: oled_colour = 16'b00011_001000_00101; 
		3353: oled_colour = 16'b00010_001000_00110; 
		3354: oled_colour = 16'b00111_010001_01010; 
		3355: oled_colour = 16'b10000_100000_01110; 
		3356: oled_colour = 16'b01111_011111_01110; 
		3357: oled_colour = 16'b10000_100010_01111; 
		3358: oled_colour = 16'b10000_100001_01110; 
		3359: oled_colour = 16'b01111_011111_01110; 
		3360: oled_colour = 16'b00011_001000_00110; 
		3361: oled_colour = 16'b00100_001000_00101; 
		3362: oled_colour = 16'b01100_011010_01110; 
		3363: oled_colour = 16'b00110_001101_01000; 
		3364: oled_colour = 16'b00100_001010_00111; 
		3365: oled_colour = 16'b00011_000101_00011; 
		3366: oled_colour = 16'b00011_000101_00011; 
		3367: oled_colour = 16'b00011_000101_00011; 
		3368: oled_colour = 16'b00011_000101_00011; 
		3369: oled_colour = 16'b00011_000101_00011; 
		3370: oled_colour = 16'b00011_000101_00010; 
		3371: oled_colour = 16'b00011_000101_00011; 
		3372: oled_colour = 16'b00010_000100_00011; 
		3373: oled_colour = 16'b00010_000100_00011; 
		3374: oled_colour = 16'b00011_000111_00101; 
		3375: oled_colour = 16'b00111_001101_00111; 
		3376: oled_colour = 16'b01010_010011_01000; 
		3377: oled_colour = 16'b01001_010010_00111; 
		3378: oled_colour = 16'b01000_001111_00110; 
		3379: oled_colour = 16'b00100_001000_00100; 
		3380: oled_colour = 16'b00001_000001_00010; 
		3381: oled_colour = 16'b00101_001011_00111; 
		3382: oled_colour = 16'b00110_001110_01001; 
		3383: oled_colour = 16'b01101_011011_01101; 
		3384: oled_colour = 16'b11010_110100_10011; 
		3385: oled_colour = 16'b11100_110110_10011; 
		3386: oled_colour = 16'b11000_101111_10001; 
		3387: oled_colour = 16'b10010_100101_10000; 
		3388: oled_colour = 16'b10000_100001_10000; 
		3389: oled_colour = 16'b01101_011010_01110; 
		3390: oled_colour = 16'b01011_011000_01100; 
		3391: oled_colour = 16'b01100_011001_01101; 
		3392: oled_colour = 16'b01100_011001_01101; 
		3393: oled_colour = 16'b01100_011001_01101; 
		3394: oled_colour = 16'b01100_011000_01100; 
		3395: oled_colour = 16'b01100_011001_01100; 
		3396: oled_colour = 16'b01100_011001_01101; 
		3397: oled_colour = 16'b01100_011000_01101; 
		3398: oled_colour = 16'b01100_011000_01100; 
		3399: oled_colour = 16'b01100_011000_01100; 
		3400: oled_colour = 16'b01100_011000_01101; 
		3401: oled_colour = 16'b01100_011000_01101; 
		3402: oled_colour = 16'b01100_011000_01101; 
		3403: oled_colour = 16'b01100_011000_01101; 
		3404: oled_colour = 16'b01011_011000_01101; 
		3405: oled_colour = 16'b01100_011001_01101; 
		3406: oled_colour = 16'b01101_011010_01110; 
		3407: oled_colour = 16'b01101_011010_01110; 
		3408: oled_colour = 16'b01101_011010_01110; 
		3409: oled_colour = 16'b01101_011011_01110; 
		3410: oled_colour = 16'b01101_011010_01110; 
		3411: oled_colour = 16'b01101_011011_01110; 
		3412: oled_colour = 16'b01101_011011_01110; 
		3413: oled_colour = 16'b01101_011010_01110; 
		3414: oled_colour = 16'b01101_011010_01101; 
		3415: oled_colour = 16'b01101_011010_01101; 
		3416: oled_colour = 16'b01101_011010_01101; 
		3417: oled_colour = 16'b01101_011010_01101; 
		3418: oled_colour = 16'b01101_011010_01101; 
		3419: oled_colour = 16'b01101_011010_01101; 
		3420: oled_colour = 16'b01101_011010_01101; 
		3421: oled_colour = 16'b01101_011010_01110; 
		3422: oled_colour = 16'b01101_011010_01110; 
		3423: oled_colour = 16'b01101_011010_01101; 
		3424: oled_colour = 16'b01101_011010_01101; 
		3425: oled_colour = 16'b01101_011001_01101; 
		3426: oled_colour = 16'b01101_011010_01110; 
		3427: oled_colour = 16'b01101_011011_01110; 
		3428: oled_colour = 16'b01100_011010_01101; 
		3429: oled_colour = 16'b01101_011010_01110; 
		3430: oled_colour = 16'b01101_011010_01110; 
		3431: oled_colour = 16'b01100_011000_01100; 
		3432: oled_colour = 16'b01100_011000_01101; 
		3433: oled_colour = 16'b01100_011000_01101; 
		3434: oled_colour = 16'b01100_011001_01101; 
		3435: oled_colour = 16'b01100_011000_01101; 
		3436: oled_colour = 16'b01100_011000_01101; 
		3437: oled_colour = 16'b01100_011001_01101; 
		3438: oled_colour = 16'b01101_011010_01110; 
		3439: oled_colour = 16'b01101_011011_01110; 
		3440: oled_colour = 16'b01101_011011_01110; 
		3441: oled_colour = 16'b01101_011010_01110; 
		3442: oled_colour = 16'b01101_011011_01110; 
		3443: oled_colour = 16'b01110_011100_01110; 
		3444: oled_colour = 16'b01000_010001_01010; 
		3445: oled_colour = 16'b00101_001100_01001; 
		3446: oled_colour = 16'b00100_001101_01001; 
		3447: oled_colour = 16'b00100_001011_01000; 
		3448: oled_colour = 16'b00011_001001_00110; 
		3449: oled_colour = 16'b00010_001000_00101; 
		3450: oled_colour = 16'b00101_001110_01001; 
		3451: oled_colour = 16'b01110_011101_01110; 
		3452: oled_colour = 16'b01101_011010_01100; 
		3453: oled_colour = 16'b01100_011001_01100; 
		3454: oled_colour = 16'b01101_011011_01100; 
		3455: oled_colour = 16'b01011_011000_01011; 
		3456: oled_colour = 16'b00100_001001_00101; 
		3457: oled_colour = 16'b00100_001000_00110; 
		3458: oled_colour = 16'b00100_001010_00111; 
		3459: oled_colour = 16'b00100_001010_00111; 
		3460: oled_colour = 16'b00101_001110_01001; 
		3461: oled_colour = 16'b00010_000101_00011; 
		3462: oled_colour = 16'b00010_000011_00010; 
		3463: oled_colour = 16'b00011_000100_00010; 
		3464: oled_colour = 16'b00011_000101_00011; 
		3465: oled_colour = 16'b00011_000101_00011; 
		3466: oled_colour = 16'b00011_000101_00011; 
		3467: oled_colour = 16'b00011_000101_00011; 
		3468: oled_colour = 16'b00010_000100_00010; 
		3469: oled_colour = 16'b00101_001010_00110; 
		3470: oled_colour = 16'b01000_010001_01001; 
		3471: oled_colour = 16'b00111_001111_00111; 
		3472: oled_colour = 16'b01000_010010_01000; 
		3473: oled_colour = 16'b01010_010110_01010; 
		3474: oled_colour = 16'b00110_001101_00111; 
		3475: oled_colour = 16'b01001_010010_01000; 
		3476: oled_colour = 16'b00111_001101_00111; 
		3477: oled_colour = 16'b00010_000100_00011; 
		3478: oled_colour = 16'b00010_000100_00011; 
		3479: oled_colour = 16'b00100_001010_00111; 
		3480: oled_colour = 16'b01010_010110_01100; 
		3481: oled_colour = 16'b10011_100111_10000; 
		3482: oled_colour = 16'b11001_110010_10010; 
		3483: oled_colour = 16'b11101_111000_10100; 
		3484: oled_colour = 16'b10101_101001_10000; 
		3485: oled_colour = 16'b00101_001101_01000; 
		3486: oled_colour = 16'b00111_010001_01010; 
		3487: oled_colour = 16'b00100_001011_01000; 
		3488: oled_colour = 16'b00101_001101_01001; 
		3489: oled_colour = 16'b00101_001110_01001; 
		3490: oled_colour = 16'b00100_001100_01000; 
		3491: oled_colour = 16'b00101_001101_01000; 
		3492: oled_colour = 16'b00101_001100_01000; 
		3493: oled_colour = 16'b00101_001101_01001; 
		3494: oled_colour = 16'b00110_001111_01001; 
		3495: oled_colour = 16'b00101_001101_01000; 
		3496: oled_colour = 16'b00101_001101_01000; 
		3497: oled_colour = 16'b00110_001110_01001; 
		3498: oled_colour = 16'b00101_001110_01001; 
		3499: oled_colour = 16'b00101_001101_01000; 
		3500: oled_colour = 16'b00101_001101_01001; 
		3501: oled_colour = 16'b00110_001110_01001; 
		3502: oled_colour = 16'b00101_001101_01000; 
		3503: oled_colour = 16'b00101_001101_01000; 
		3504: oled_colour = 16'b00101_001101_01000; 
		3505: oled_colour = 16'b00101_001100_01000; 
		3506: oled_colour = 16'b00101_001101_01001; 
		3507: oled_colour = 16'b00101_001101_01001; 
		3508: oled_colour = 16'b00100_001100_01000; 
		3509: oled_colour = 16'b00101_001101_01001; 
		3510: oled_colour = 16'b00110_001110_01001; 
		3511: oled_colour = 16'b00101_001101_01001; 
		3512: oled_colour = 16'b00100_001100_01000; 
		3513: oled_colour = 16'b00101_001110_01001; 
		3514: oled_colour = 16'b00101_001110_01001; 
		3515: oled_colour = 16'b00101_001100_01000; 
		3516: oled_colour = 16'b00101_001101_01000; 
		3517: oled_colour = 16'b00101_001100_01000; 
		3518: oled_colour = 16'b00101_001101_01001; 
		3519: oled_colour = 16'b00110_001110_01001; 
		3520: oled_colour = 16'b00101_001101_01000; 
		3521: oled_colour = 16'b00101_001101_01000; 
		3522: oled_colour = 16'b00101_001101_01000; 
		3523: oled_colour = 16'b00101_001110_01001; 
		3524: oled_colour = 16'b00100_001100_01000; 
		3525: oled_colour = 16'b00101_001101_01000; 
		3526: oled_colour = 16'b00110_001110_01001; 
		3527: oled_colour = 16'b00101_001101_01000; 
		3528: oled_colour = 16'b00101_001101_01000; 
		3529: oled_colour = 16'b00101_001101_01000; 
		3530: oled_colour = 16'b00101_001100_01000; 
		3531: oled_colour = 16'b00101_001110_01001; 
		3532: oled_colour = 16'b00110_001110_01001; 
		3533: oled_colour = 16'b00101_001101_01000; 
		3534: oled_colour = 16'b00101_001101_01000; 
		3535: oled_colour = 16'b00101_001110_01000; 
		3536: oled_colour = 16'b00101_001101_01001; 
		3537: oled_colour = 16'b00100_001100_01000; 
		3538: oled_colour = 16'b00101_001101_01001; 
		3539: oled_colour = 16'b00101_001101_01001; 
		3540: oled_colour = 16'b00011_001011_00111; 
		3541: oled_colour = 16'b00011_001010_00111; 
		3542: oled_colour = 16'b00011_001010_00111; 
		3543: oled_colour = 16'b00100_001011_00111; 
		3544: oled_colour = 16'b00100_001011_00111; 
		3545: oled_colour = 16'b00011_001000_00101; 
		3546: oled_colour = 16'b00010_001001_00111; 
		3547: oled_colour = 16'b01101_011100_01110; 
		3548: oled_colour = 16'b10100_101000_10000; 
		3549: oled_colour = 16'b10100_100111_10000; 
		3550: oled_colour = 16'b10100_100111_10000; 
		3551: oled_colour = 16'b10001_100010_01111; 
		3552: oled_colour = 16'b01000_010100_01011; 
		3553: oled_colour = 16'b00110_001110_01000; 
		3554: oled_colour = 16'b00010_000011_00011; 
		3555: oled_colour = 16'b00101_001011_00111; 
		3556: oled_colour = 16'b01111_100001_01111; 
		3557: oled_colour = 16'b01101_011101_01101; 
		3558: oled_colour = 16'b00110_001101_00111; 
		3559: oled_colour = 16'b00011_000110_00100; 
		3560: oled_colour = 16'b00010_000100_00010; 
		3561: oled_colour = 16'b00010_000100_00010; 
		3562: oled_colour = 16'b00011_000101_00011; 
		3563: oled_colour = 16'b00010_000100_00010; 
		3564: oled_colour = 16'b00100_001000_00101; 
		3565: oled_colour = 16'b00100_001011_00111; 
		3566: oled_colour = 16'b00111_010001_01001; 
		3567: oled_colour = 16'b01001_010100_01011; 
		3568: oled_colour = 16'b00110_001111_01010; 
		3569: oled_colour = 16'b01000_010100_01100; 
		3570: oled_colour = 16'b00101_001110_01001; 
		3571: oled_colour = 16'b01000_010011_01010; 
		3572: oled_colour = 16'b00101_001100_00111; 
		3573: oled_colour = 16'b00100_001010_00110; 
		3574: oled_colour = 16'b00010_000101_00011; 
		3575: oled_colour = 16'b00010_000100_00010; 
		3576: oled_colour = 16'b00010_000101_00100; 
		3577: oled_colour = 16'b00100_001010_00111; 
		3578: oled_colour = 16'b01001_010100_01011; 
		3579: oled_colour = 16'b10011_100111_10000; 
		3580: oled_colour = 16'b01110_011110_01101; 
		3581: oled_colour = 16'b01111_011111_01110; 
		3582: oled_colour = 16'b11001_110001_10011; 
		3583: oled_colour = 16'b10000_100010_01111; 
		3584: oled_colour = 16'b01011_011001_01101; 
		3585: oled_colour = 16'b01000_010011_01011; 
		3586: oled_colour = 16'b00101_001111_01001; 
		3587: oled_colour = 16'b00101_001111_01001; 
		3588: oled_colour = 16'b01010_010110_01011; 
		3589: oled_colour = 16'b00110_001111_01001; 
		3590: oled_colour = 16'b00101_001110_01000; 
		3591: oled_colour = 16'b01000_010011_01010; 
		3592: oled_colour = 16'b00110_010000_01001; 
		3593: oled_colour = 16'b00100_001101_01000; 
		3594: oled_colour = 16'b01000_010011_01010; 
		3595: oled_colour = 16'b00111_010001_01001; 
		3596: oled_colour = 16'b00100_001101_01000; 
		3597: oled_colour = 16'b00111_010010_01010; 
		3598: oled_colour = 16'b00111_010010_01010; 
		3599: oled_colour = 16'b00100_001101_01000; 
		3600: oled_colour = 16'b00111_010010_01010; 
		3601: oled_colour = 16'b01000_010100_01010; 
		3602: oled_colour = 16'b00100_001101_01000; 
		3603: oled_colour = 16'b00111_010000_01001; 
		3604: oled_colour = 16'b01000_010011_01010; 
		3605: oled_colour = 16'b00101_001110_01000; 
		3606: oled_colour = 16'b00110_010000_01001; 
		3607: oled_colour = 16'b01001_010100_01011; 
		3608: oled_colour = 16'b00101_001110_01000; 
		3609: oled_colour = 16'b00101_001111_01001; 
		3610: oled_colour = 16'b01000_010011_01010; 
		3611: oled_colour = 16'b00101_001111_01001; 
		3612: oled_colour = 16'b00101_001110_01001; 
		3613: oled_colour = 16'b01001_010101_01011; 
		3614: oled_colour = 16'b00110_001111_01001; 
		3615: oled_colour = 16'b00101_001110_01000; 
		3616: oled_colour = 16'b01000_010011_01010; 
		3617: oled_colour = 16'b00110_010000_01001; 
		3618: oled_colour = 16'b00101_001110_01000; 
		3619: oled_colour = 16'b01000_010011_01010; 
		3620: oled_colour = 16'b00111_010001_01001; 
		3621: oled_colour = 16'b00100_001101_01001; 
		3622: oled_colour = 16'b01000_010010_01010; 
		3623: oled_colour = 16'b00111_010010_01010; 
		3624: oled_colour = 16'b00100_001101_01000; 
		3625: oled_colour = 16'b01000_010011_01010; 
		3626: oled_colour = 16'b01001_010100_01011; 
		3627: oled_colour = 16'b00100_001101_01000; 
		3628: oled_colour = 16'b00111_010001_01001; 
		3629: oled_colour = 16'b01000_010011_01010; 
		3630: oled_colour = 16'b00101_001110_01000; 
		3631: oled_colour = 16'b00110_010000_01001; 
		3632: oled_colour = 16'b01001_010100_01011; 
		3633: oled_colour = 16'b00101_001110_01000; 
		3634: oled_colour = 16'b00101_001111_01001; 
		3635: oled_colour = 16'b01000_010100_01011; 
		3636: oled_colour = 16'b00100_001100_01000; 
		3637: oled_colour = 16'b00011_001001_00111; 
		3638: oled_colour = 16'b00101_001101_01000; 
		3639: oled_colour = 16'b00011_001010_00111; 
		3640: oled_colour = 16'b00011_001000_00110; 
		3641: oled_colour = 16'b00011_000111_00101; 
		3642: oled_colour = 16'b00011_001000_00101; 
		3643: oled_colour = 16'b00111_010001_01010; 
		3644: oled_colour = 16'b01101_011010_01101; 
		3645: oled_colour = 16'b01100_011001_01100; 
		3646: oled_colour = 16'b01101_011010_01101; 
		3647: oled_colour = 16'b01110_011100_01101; 
		3648: oled_colour = 16'b00011_000111_00101; 
		3649: oled_colour = 16'b00011_001001_00110; 
		3650: oled_colour = 16'b00101_001100_01000; 
		3651: oled_colour = 16'b00011_000111_00110; 
		3652: oled_colour = 16'b00111_001111_01000; 
		3653: oled_colour = 16'b10110_101101_10010; 
		3654: oled_colour = 16'b10011_101000_10000; 
		3655: oled_colour = 16'b01011_011001_01100; 
		3656: oled_colour = 16'b00110_001101_01000; 
		3657: oled_colour = 16'b00011_000110_00100; 
		3658: oled_colour = 16'b00001_000011_00010; 
		3659: oled_colour = 16'b00011_000110_00100; 
		3660: oled_colour = 16'b00101_001101_01000; 
		3661: oled_colour = 16'b00101_001101_01000; 
		3662: oled_colour = 16'b00101_001011_01000; 
		3663: oled_colour = 16'b00110_001110_01001; 
		3664: oled_colour = 16'b00011_000111_00101; 
		3665: oled_colour = 16'b00011_000110_00101; 
		3666: oled_colour = 16'b00100_001010_00111; 
		3667: oled_colour = 16'b00101_001011_01000; 
		3668: oled_colour = 16'b00100_001010_00110; 
		3669: oled_colour = 16'b00101_001110_01000; 
		3670: oled_colour = 16'b00100_001001_00110; 
		3671: oled_colour = 16'b00011_000101_00100; 
		3672: oled_colour = 16'b00011_000101_00010; 
		3673: oled_colour = 16'b00010_000100_00010; 
		3674: oled_colour = 16'b00010_000100_00011; 
		3675: oled_colour = 16'b00011_001001_00111; 
		3676: oled_colour = 16'b00011_001001_00111; 
		3677: oled_colour = 16'b01010_011000_01100; 
		3678: oled_colour = 16'b10110_101101_10010; 
		3679: oled_colour = 16'b11100_110111_10100; 
		3680: oled_colour = 16'b11001_110001_10010; 
		3681: oled_colour = 16'b10011_100110_10000; 
		3682: oled_colour = 16'b01100_011100_01101; 
		3683: oled_colour = 16'b00100_001100_01000; 
		3684: oled_colour = 16'b10000_100010_01110; 
		3685: oled_colour = 16'b01000_010010_01010; 
		3686: oled_colour = 16'b00100_001011_01000; 
		3687: oled_colour = 16'b01111_011111_01110; 
		3688: oled_colour = 16'b01001_010101_01010; 
		3689: oled_colour = 16'b00011_001001_01000; 
		3690: oled_colour = 16'b01110_011110_01110; 
		3691: oled_colour = 16'b01100_011001_01100; 
		3692: oled_colour = 16'b00011_001001_00111; 
		3693: oled_colour = 16'b01100_011010_01100; 
		3694: oled_colour = 16'b01100_011001_01100; 
		3695: oled_colour = 16'b00011_001001_00111; 
		3696: oled_colour = 16'b01010_010111_01100; 
		3697: oled_colour = 16'b01111_011111_01110; 
		3698: oled_colour = 16'b00011_001010_00111; 
		3699: oled_colour = 16'b01001_010100_01011; 
		3700: oled_colour = 16'b01111_100000_01110; 
		3701: oled_colour = 16'b00100_001011_01000; 
		3702: oled_colour = 16'b00111_010001_01010; 
		3703: oled_colour = 16'b10000_100001_01111; 
		3704: oled_colour = 16'b00101_001101_01001; 
		3705: oled_colour = 16'b00110_001111_01001; 
		3706: oled_colour = 16'b01111_011111_01110; 
		3707: oled_colour = 16'b00110_001110_01001; 
		3708: oled_colour = 16'b00101_001101_01001; 
		3709: oled_colour = 16'b10000_100001_01111; 
		3710: oled_colour = 16'b00111_010001_01010; 
		3711: oled_colour = 16'b00100_001100_01000; 
		3712: oled_colour = 16'b01111_011111_01110; 
		3713: oled_colour = 16'b01001_010100_01011; 
		3714: oled_colour = 16'b00011_001001_00111; 
		3715: oled_colour = 16'b01111_011110_01110; 
		3716: oled_colour = 16'b01011_011000_01011; 
		3717: oled_colour = 16'b00011_001001_00111; 
		3718: oled_colour = 16'b01100_011010_01101; 
		3719: oled_colour = 16'b01011_011001_01100; 
		3720: oled_colour = 16'b00011_001001_00111; 
		3721: oled_colour = 16'b01011_011000_01100; 
		3722: oled_colour = 16'b01111_011111_01110; 
		3723: oled_colour = 16'b00011_001010_01000; 
		3724: oled_colour = 16'b01001_010101_01011; 
		3725: oled_colour = 16'b01111_100000_01110; 
		3726: oled_colour = 16'b00100_001011_01000; 
		3727: oled_colour = 16'b00111_010001_01010; 
		3728: oled_colour = 16'b10001_100010_01111; 
		3729: oled_colour = 16'b00101_001101_01000; 
		3730: oled_colour = 16'b00110_001110_01001; 
		3731: oled_colour = 16'b01111_100000_01110; 
		3732: oled_colour = 16'b00110_001110_01001; 
		3733: oled_colour = 16'b00010_001000_00110; 
		3734: oled_colour = 16'b00111_010001_01010; 
		3735: oled_colour = 16'b00100_001011_01000; 
		3736: oled_colour = 16'b00010_001000_00110; 
		3737: oled_colour = 16'b00100_001011_00111; 
		3738: oled_colour = 16'b00011_001001_00110; 
		3739: oled_colour = 16'b00011_001010_00111; 
		3740: oled_colour = 16'b01111_011111_01110; 
		3741: oled_colour = 16'b10110_101011_10001; 
		3742: oled_colour = 16'b10101_101001_10000; 
		3743: oled_colour = 16'b10100_100110_01111; 
		3744: oled_colour = 16'b00100_001010_00111; 
		3745: oled_colour = 16'b00100_001011_00111; 
		3746: oled_colour = 16'b00011_000110_00101; 
		3747: oled_colour = 16'b01000_010010_01010; 
		3748: oled_colour = 16'b00110_010000_01010; 
		3749: oled_colour = 16'b00101_001100_01000; 
		3750: oled_colour = 16'b10010_100110_01111; 
		3751: oled_colour = 16'b11000_110000_10010; 
		3752: oled_colour = 16'b10010_100101_10000; 
		3753: oled_colour = 16'b01110_011101_01101; 
		3754: oled_colour = 16'b01010_010110_01010; 
		3755: oled_colour = 16'b00101_001100_01000; 
		3756: oled_colour = 16'b00101_001101_01000; 
		3757: oled_colour = 16'b01000_010100_01011; 
		3758: oled_colour = 16'b00011_001000_00110; 
		3759: oled_colour = 16'b00110_001110_01000; 
		3760: oled_colour = 16'b01001_010011_01010; 
		3761: oled_colour = 16'b00110_001101_00111; 
		3762: oled_colour = 16'b00100_001010_00111; 
		3763: oled_colour = 16'b00011_001001_00110; 
		3764: oled_colour = 16'b00111_010010_01010; 
		3765: oled_colour = 16'b01001_010110_01100; 
		3766: oled_colour = 16'b00100_001011_01000; 
		3767: oled_colour = 16'b00011_001000_00110; 
		3768: oled_colour = 16'b00010_000110_00100; 
		3769: oled_colour = 16'b00011_000110_00100; 
		3770: oled_colour = 16'b00011_000101_00011; 
		3771: oled_colour = 16'b00010_000100_00010; 
		3772: oled_colour = 16'b00010_000101_00011; 
		3773: oled_colour = 16'b00011_001000_00110; 
		3774: oled_colour = 16'b00110_010000_01010; 
		3775: oled_colour = 16'b01110_011110_01110; 
		3776: oled_colour = 16'b10111_101110_10001; 
		3777: oled_colour = 16'b11110_111010_10100; 
		3778: oled_colour = 16'b10001_100001_01101; 
		3779: oled_colour = 16'b01011_011000_01011; 
		3780: oled_colour = 16'b01110_011110_01101; 
		3781: oled_colour = 16'b01000_010010_01011; 
		3782: oled_colour = 16'b00101_001101_01001; 
		3783: oled_colour = 16'b01110_011110_01110; 
		3784: oled_colour = 16'b01011_010111_01100; 
		3785: oled_colour = 16'b00110_001110_01001; 
		3786: oled_colour = 16'b01100_011010_01100; 
		3787: oled_colour = 16'b01011_011000_01100; 
		3788: oled_colour = 16'b00110_001110_01001; 
		3789: oled_colour = 16'b01110_011101_01101; 
		3790: oled_colour = 16'b01110_011100_01101; 
		3791: oled_colour = 16'b00110_001110_01010; 
		3792: oled_colour = 16'b01010_010101_01011; 
		3793: oled_colour = 16'b01100_011001_01100; 
		3794: oled_colour = 16'b00111_001111_01010; 
		3795: oled_colour = 16'b01001_010100_01011; 
		3796: oled_colour = 16'b01111_011110_01110; 
		3797: oled_colour = 16'b00111_001111_01010; 
		3798: oled_colour = 16'b01000_010010_01010; 
		3799: oled_colour = 16'b01101_011100_01101; 
		3800: oled_colour = 16'b00111_010000_01010; 
		3801: oled_colour = 16'b01000_010010_01011; 
		3802: oled_colour = 16'b10000_100001_01111; 
		3803: oled_colour = 16'b01001_010010_01011; 
		3804: oled_colour = 16'b00111_010000_01010; 
		3805: oled_colour = 16'b01100_011010_01100; 
		3806: oled_colour = 16'b01001_010011_01011; 
		3807: oled_colour = 16'b00111_001111_01010; 
		3808: oled_colour = 16'b01110_011101_01101; 
		3809: oled_colour = 16'b01010_010110_01100; 
		3810: oled_colour = 16'b00110_001110_01001; 
		3811: oled_colour = 16'b01101_011010_01100; 
		3812: oled_colour = 16'b01011_011000_01100; 
		3813: oled_colour = 16'b00110_001101_01001; 
		3814: oled_colour = 16'b01111_011101_01101; 
		3815: oled_colour = 16'b01101_011011_01101; 
		3816: oled_colour = 16'b00110_001110_01010; 
		3817: oled_colour = 16'b01010_010110_01011; 
		3818: oled_colour = 16'b01100_011001_01100; 
		3819: oled_colour = 16'b00110_001111_01010; 
		3820: oled_colour = 16'b01010_010101_01011; 
		3821: oled_colour = 16'b01111_011111_01110; 
		3822: oled_colour = 16'b00111_001111_01010; 
		3823: oled_colour = 16'b01000_010010_01010; 
		3824: oled_colour = 16'b01110_011101_01101; 
		3825: oled_colour = 16'b01000_010001_01010; 
		3826: oled_colour = 16'b01000_010010_01010; 
		3827: oled_colour = 16'b10010_100011_01111; 
		3828: oled_colour = 16'b01001_010010_01010; 
		3829: oled_colour = 16'b00011_001011_00111; 
		3830: oled_colour = 16'b00101_001101_01000; 
		3831: oled_colour = 16'b00100_001101_01000; 
		3832: oled_colour = 16'b00011_001010_00111; 
		3833: oled_colour = 16'b00100_001010_00111; 
		3834: oled_colour = 16'b00011_001001_00111; 
		3835: oled_colour = 16'b00011_001010_00111; 
		3836: oled_colour = 16'b01000_010001_01010; 
		3837: oled_colour = 16'b01101_011011_01101; 
		3838: oled_colour = 16'b01101_011011_01100; 
		3839: oled_colour = 16'b10000_100000_01110; 
		3840: oled_colour = 16'b00011_001000_00101; 
		3841: oled_colour = 16'b00011_000101_00011; 
		3842: oled_colour = 16'b00001_000001_00010; 
		3843: oled_colour = 16'b01101_011100_01101; 
		3844: oled_colour = 16'b10101_101011_10001; 
		3845: oled_colour = 16'b01000_010011_01011; 
		3846: oled_colour = 16'b00101_001101_01001; 
		3847: oled_colour = 16'b01010_010101_01010; 
		3848: oled_colour = 16'b01111_011110_01101; 
		3849: oled_colour = 16'b10011_100110_01111; 
		3850: oled_colour = 16'b10100_101000_10000; 
		3851: oled_colour = 16'b00110_001101_01000; 
		3852: oled_colour = 16'b00010_000101_00101; 
		3853: oled_colour = 16'b00011_000111_00101; 
		3854: oled_colour = 16'b00101_001010_00110; 
		3855: oled_colour = 16'b00111_010001_01011; 
		3856: oled_colour = 16'b00110_010000_01010; 
		3857: oled_colour = 16'b00100_001101_01001; 
		3858: oled_colour = 16'b00011_001001_00111; 
		3859: oled_colour = 16'b00101_001110_01001; 
		3860: oled_colour = 16'b00100_001010_01000; 
		3861: oled_colour = 16'b00011_001001_00111; 
		3862: oled_colour = 16'b00011_001000_00110; 
		3863: oled_colour = 16'b00011_001000_00110; 
		3864: oled_colour = 16'b00010_000100_00100; 
		3865: oled_colour = 16'b00011_000110_00101; 
		3866: oled_colour = 16'b00011_000110_00100; 
		3867: oled_colour = 16'b00011_000110_00100; 
		3868: oled_colour = 16'b00011_000101_00011; 
		3869: oled_colour = 16'b00010_000100_00010; 
		3870: oled_colour = 16'b00010_000101_00011; 
		3871: oled_colour = 16'b00011_001000_00110; 
		3872: oled_colour = 16'b00111_010001_01010; 
		3873: oled_colour = 16'b10001_100011_01111; 
		3874: oled_colour = 16'b01001_010101_01010; 
		3875: oled_colour = 16'b10111_101110_10010; 
		3876: oled_colour = 16'b11010_110011_10011; 
		3877: oled_colour = 16'b10011_100110_10000; 
		3878: oled_colour = 16'b01100_011001_01101; 
		3879: oled_colour = 16'b10000_100000_01111; 
		3880: oled_colour = 16'b01010_010111_01100; 
		3881: oled_colour = 16'b00101_001101_01001; 
		3882: oled_colour = 16'b01110_011100_01101; 
		3883: oled_colour = 16'b01100_011001_01100; 
		3884: oled_colour = 16'b00101_001110_01001; 
		3885: oled_colour = 16'b01010_010110_01011; 
		3886: oled_colour = 16'b01011_010110_01100; 
		3887: oled_colour = 16'b00110_001110_01001; 
		3888: oled_colour = 16'b01011_010110_01011; 
		3889: oled_colour = 16'b01101_011011_01101; 
		3890: oled_colour = 16'b00101_001101_01001; 
		3891: oled_colour = 16'b01010_010101_01011; 
		3892: oled_colour = 16'b10001_100010_01111; 
		3893: oled_colour = 16'b00111_001111_01010; 
		3894: oled_colour = 16'b01000_010010_01010; 
		3895: oled_colour = 16'b01111_011110_01110; 
		3896: oled_colour = 16'b00111_010000_01001; 
		3897: oled_colour = 16'b00111_010001_01010; 
		3898: oled_colour = 16'b01100_011000_01101; 
		3899: oled_colour = 16'b01000_010001_01010; 
		3900: oled_colour = 16'b00111_001111_01001; 
		3901: oled_colour = 16'b01110_011101_01101; 
		3902: oled_colour = 16'b01001_010010_01010; 
		3903: oled_colour = 16'b00110_001101_01001; 
		3904: oled_colour = 16'b10000_100000_01110; 
		3905: oled_colour = 16'b01011_010111_01100; 
		3906: oled_colour = 16'b00101_001101_01001; 
		3907: oled_colour = 16'b01110_011100_01101; 
		3908: oled_colour = 16'b01011_011000_01011; 
		3909: oled_colour = 16'b00110_001101_01001; 
		3910: oled_colour = 16'b01010_010110_01100; 
		3911: oled_colour = 16'b01010_010110_01100; 
		3912: oled_colour = 16'b00110_001110_01001; 
		3913: oled_colour = 16'b01011_010111_01100; 
		3914: oled_colour = 16'b01101_011011_01101; 
		3915: oled_colour = 16'b00101_001101_01001; 
		3916: oled_colour = 16'b01010_010110_01011; 
		3917: oled_colour = 16'b10010_100011_01111; 
		3918: oled_colour = 16'b00111_001110_01010; 
		3919: oled_colour = 16'b01000_010010_01010; 
		3920: oled_colour = 16'b01111_011111_01101; 
		3921: oled_colour = 16'b00111_010000_01010; 
		3922: oled_colour = 16'b00111_010000_01010; 
		3923: oled_colour = 16'b01101_011010_01101; 
		3924: oled_colour = 16'b01000_010001_01010; 
		3925: oled_colour = 16'b00011_001010_00111; 
		3926: oled_colour = 16'b00101_001110_01001; 
		3927: oled_colour = 16'b00100_001101_01000; 
		3928: oled_colour = 16'b00011_001010_00111; 
		3929: oled_colour = 16'b00100_001100_00111; 
		3930: oled_colour = 16'b00011_001001_00110; 
		3931: oled_colour = 16'b00011_001001_00110; 
		3932: oled_colour = 16'b00101_001101_01000; 
		3933: oled_colour = 16'b10011_100101_10000; 
		3934: oled_colour = 16'b10110_101011_10001; 
		3935: oled_colour = 16'b10101_101001_10001; 
		3936: oled_colour = 16'b00011_000110_00100; 
		3937: oled_colour = 16'b00011_000111_00101; 
		3938: oled_colour = 16'b00011_000111_00100; 
		3939: oled_colour = 16'b00100_001000_00101; 
		3940: oled_colour = 16'b10010_100011_01111; 
		3941: oled_colour = 16'b11000_101111_10010; 
		3942: oled_colour = 16'b10000_100010_01110; 
		3943: oled_colour = 16'b00111_010001_01010; 
		3944: oled_colour = 16'b00011_001001_00111; 
		3945: oled_colour = 16'b00011_001000_00111; 
		3946: oled_colour = 16'b00101_001100_01000; 
		3947: oled_colour = 16'b00101_001100_01000; 
		3948: oled_colour = 16'b00101_001100_01000; 
		3949: oled_colour = 16'b00011_000111_00110; 
		3950: oled_colour = 16'b00101_001100_00111; 
		3951: oled_colour = 16'b00101_001100_00111; 
		3952: oled_colour = 16'b00110_001110_01001; 
		3953: oled_colour = 16'b00110_010000_01010; 
		3954: oled_colour = 16'b00111_001111_01000; 
		3955: oled_colour = 16'b00110_001110_01001; 
		3956: oled_colour = 16'b00100_001011_01000; 
		3957: oled_colour = 16'b01001_010110_01100; 
		3958: oled_colour = 16'b00110_001110_01001; 
		3959: oled_colour = 16'b00011_001000_00110; 
		3960: oled_colour = 16'b00011_000101_00010; 
		3961: oled_colour = 16'b00011_000100_00011; 
		3962: oled_colour = 16'b00011_000101_00100; 
		3963: oled_colour = 16'b00011_000110_00101; 
		3964: oled_colour = 16'b00011_000111_00101; 
		3965: oled_colour = 16'b00011_000110_00100; 
		3966: oled_colour = 16'b00011_000101_00011; 
		3967: oled_colour = 16'b00010_000100_00010; 
		3968: oled_colour = 16'b00010_000100_00011; 
		3969: oled_colour = 16'b00010_000101_00100; 
		3970: oled_colour = 16'b00011_000111_00101; 
		3971: oled_colour = 16'b01000_010001_01010; 
		3972: oled_colour = 16'b10010_100110_10000; 
		3973: oled_colour = 16'b11011_110110_10100; 
		3974: oled_colour = 16'b11100_110111_10100; 
		3975: oled_colour = 16'b10111_101110_10001; 
		3976: oled_colour = 16'b10001_100011_01111; 
		3977: oled_colour = 16'b01011_011001_01101; 
		3978: oled_colour = 16'b01110_011101_01110; 
		3979: oled_colour = 16'b01100_011001_01100; 
		3980: oled_colour = 16'b00101_001101_01001; 
		3981: oled_colour = 16'b01011_010110_01100; 
		3982: oled_colour = 16'b01100_011000_01101; 
		3983: oled_colour = 16'b00110_001101_01001; 
		3984: oled_colour = 16'b01100_011010_01100; 
		3985: oled_colour = 16'b10000_100000_01110; 
		3986: oled_colour = 16'b00110_001101_01001; 
		3987: oled_colour = 16'b01000_010011_01010; 
		3988: oled_colour = 16'b01101_011100_01101; 
		3989: oled_colour = 16'b00111_001111_01001; 
		3990: oled_colour = 16'b01000_010010_01010; 
		3991: oled_colour = 16'b10000_100001_01110; 
		3992: oled_colour = 16'b00111_010000_01010; 
		3993: oled_colour = 16'b00111_010000_01010; 
		3994: oled_colour = 16'b01100_011010_01101; 
		3995: oled_colour = 16'b01000_010001_01010; 
		3996: oled_colour = 16'b00111_001111_01001; 
		3997: oled_colour = 16'b10001_100011_01111; 
		3998: oled_colour = 16'b01001_010100_01010; 
		3999: oled_colour = 16'b00110_001110_01001; 
		4000: oled_colour = 16'b01100_011010_01100; 
		4001: oled_colour = 16'b01010_010101_01011; 
		4002: oled_colour = 16'b00110_001101_01001; 
		4003: oled_colour = 16'b01111_011111_01110; 
		4004: oled_colour = 16'b01101_011010_01100; 
		4005: oled_colour = 16'b00101_001101_01001; 
		4006: oled_colour = 16'b01010_010111_01100; 
		4007: oled_colour = 16'b01011_010111_01100; 
		4008: oled_colour = 16'b00110_001101_01001; 
		4009: oled_colour = 16'b01101_011011_01101; 
		4010: oled_colour = 16'b10000_100001_01110; 
		4011: oled_colour = 16'b00101_001101_01001; 
		4012: oled_colour = 16'b01001_010100_01010; 
		4013: oled_colour = 16'b01101_011011_01101; 
		4014: oled_colour = 16'b00111_001111_01010; 
		4015: oled_colour = 16'b01000_010010_01010; 
		4016: oled_colour = 16'b10001_100010_01111; 
		4017: oled_colour = 16'b00111_010000_01010; 
		4018: oled_colour = 16'b00111_010000_01010; 
		4019: oled_colour = 16'b01101_011010_01101; 
		4020: oled_colour = 16'b01000_010010_01010; 
		4021: oled_colour = 16'b00100_001011_01000; 
		4022: oled_colour = 16'b00111_010001_01010; 
		4023: oled_colour = 16'b00100_001101_01000; 
		4024: oled_colour = 16'b00011_001010_00110; 
		4025: oled_colour = 16'b00011_001001_00110; 
		4026: oled_colour = 16'b00011_001000_00110; 
		4027: oled_colour = 16'b00011_001000_00110; 
		4028: oled_colour = 16'b00011_001011_00111; 
		4029: oled_colour = 16'b00111_010001_01010; 
		4030: oled_colour = 16'b01001_010100_01011; 
		4031: oled_colour = 16'b01010_010100_01010; 
		4032: oled_colour = 16'b00110_001110_01000; 
		4033: oled_colour = 16'b00011_001001_00110; 
		4034: oled_colour = 16'b00100_001010_00111; 
		4035: oled_colour = 16'b00011_000101_00011; 
		4036: oled_colour = 16'b00010_000101_00100; 
		4037: oled_colour = 16'b01001_010100_01001; 
		4038: oled_colour = 16'b10010_100100_01111; 
		4039: oled_colour = 16'b10111_101101_10010; 
		4040: oled_colour = 16'b10110_101100_10010; 
		4041: oled_colour = 16'b10010_100110_10000; 
		4042: oled_colour = 16'b01101_011101_01110; 
		4043: oled_colour = 16'b00100_001011_01000; 
		4044: oled_colour = 16'b00110_001111_01001; 
		4045: oled_colour = 16'b00100_001011_00111; 
		4046: oled_colour = 16'b00101_001110_01001; 
		4047: oled_colour = 16'b01010_010111_01100; 
		4048: oled_colour = 16'b01000_010001_01010; 
		4049: oled_colour = 16'b00110_001110_01000; 
		4050: oled_colour = 16'b01011_011001_01101; 
		4051: oled_colour = 16'b00111_010010_01011; 
		4052: oled_colour = 16'b00011_000111_00101; 
		4053: oled_colour = 16'b00100_001010_00111; 
		4054: oled_colour = 16'b00100_001011_01000; 
		4055: oled_colour = 16'b00100_001010_00111; 
		4056: oled_colour = 16'b00011_000101_00011; 
		4057: oled_colour = 16'b00011_000101_00011; 
		4058: oled_colour = 16'b00011_000101_00011; 
		4059: oled_colour = 16'b00010_000101_00011; 
		4060: oled_colour = 16'b00010_000101_00011; 
		4061: oled_colour = 16'b00011_000101_00100; 
		4062: oled_colour = 16'b00011_000110_00101; 
		4063: oled_colour = 16'b00011_000111_00101; 
		4064: oled_colour = 16'b00011_000101_00011; 
		4065: oled_colour = 16'b00011_000101_00010; 
		4066: oled_colour = 16'b00011_000101_00010; 
		4067: oled_colour = 16'b00001_000011_00010; 
		4068: oled_colour = 16'b00010_000110_00101; 
		4069: oled_colour = 16'b01001_010100_01010; 
		4070: oled_colour = 16'b10011_100111_10000; 
		4071: oled_colour = 16'b11010_110100_10011; 
		4072: oled_colour = 16'b11110_111010_10100; 
		4073: oled_colour = 16'b10010_100101_01111; 
		4074: oled_colour = 16'b01011_010111_01011; 
		4075: oled_colour = 16'b01100_011010_01101; 
		4076: oled_colour = 16'b00101_001101_01001; 
		4077: oled_colour = 16'b01001_010100_01011; 
		4078: oled_colour = 16'b01011_010110_01100; 
		4079: oled_colour = 16'b00110_001101_01001; 
		4080: oled_colour = 16'b01010_010101_01011; 
		4081: oled_colour = 16'b01101_011010_01100; 
		4082: oled_colour = 16'b00110_001110_01001; 
		4083: oled_colour = 16'b01000_010011_01010; 
		4084: oled_colour = 16'b01101_011011_01101; 
		4085: oled_colour = 16'b00110_001111_01001; 
		4086: oled_colour = 16'b01000_010010_01010; 
		4087: oled_colour = 16'b01110_011110_01110; 
		4088: oled_colour = 16'b00111_010000_01001; 
		4089: oled_colour = 16'b00111_010000_01010; 
		4090: oled_colour = 16'b01011_010111_01100; 
		4091: oled_colour = 16'b01000_010001_01010; 
		4092: oled_colour = 16'b00110_001111_01001; 
		4093: oled_colour = 16'b01101_011100_01101; 
		4094: oled_colour = 16'b01001_010011_01010; 
		4095: oled_colour = 16'b00110_001110_01001; 
		4096: oled_colour = 16'b01101_011010_01101; 
		4097: oled_colour = 16'b01001_010100_01011; 
		4098: oled_colour = 16'b00110_001101_01001; 
		4099: oled_colour = 16'b01110_011100_01101; 
		4100: oled_colour = 16'b01011_011000_01100; 
		4101: oled_colour = 16'b00110_001101_01001; 
		4102: oled_colour = 16'b01010_010101_01011; 
		4103: oled_colour = 16'b01010_010110_01011; 
		4104: oled_colour = 16'b00110_001110_01001; 
		4105: oled_colour = 16'b01010_010110_01011; 
		4106: oled_colour = 16'b01101_011010_01100; 
		4107: oled_colour = 16'b00110_001110_01001; 
		4108: oled_colour = 16'b01001_010100_01011; 
		4109: oled_colour = 16'b01101_011100_01101; 
		4110: oled_colour = 16'b00110_001111_01001; 
		4111: oled_colour = 16'b01000_010010_01010; 
		4112: oled_colour = 16'b01111_011111_01110; 
		4113: oled_colour = 16'b00111_010000_01010; 
		4114: oled_colour = 16'b00111_010000_01001; 
		4115: oled_colour = 16'b01100_011000_01100; 
		4116: oled_colour = 16'b01000_010010_01010; 
		4117: oled_colour = 16'b00100_001100_01000; 
		4118: oled_colour = 16'b00101_001101_01000; 
		4119: oled_colour = 16'b00100_001101_01000; 
		4120: oled_colour = 16'b00011_001010_00111; 
		4121: oled_colour = 16'b00011_001001_00110; 
		4122: oled_colour = 16'b00011_000111_00101; 
		4123: oled_colour = 16'b00011_000110_00100; 
		4124: oled_colour = 16'b00011_001001_00110; 
		4125: oled_colour = 16'b00101_001110_01001; 
		4126: oled_colour = 16'b10101_101001_10001; 
		4127: oled_colour = 16'b11001_110000_10010; 
		4128: oled_colour = 16'b00100_001010_00110; 
		4129: oled_colour = 16'b00101_001101_01000; 
		4130: oled_colour = 16'b00011_001000_00101; 
		4131: oled_colour = 16'b00100_001001_00110; 
		4132: oled_colour = 16'b00100_001001_00110; 
		4133: oled_colour = 16'b00001_000011_00010; 
		4134: oled_colour = 16'b00010_000101_00100; 
		4135: oled_colour = 16'b00110_001101_00111; 
		4136: oled_colour = 16'b01011_010111_01010; 
		4137: oled_colour = 16'b01111_011101_01100; 
		4138: oled_colour = 16'b01011_011000_01011; 
		4139: oled_colour = 16'b00011_001001_00111; 
		4140: oled_colour = 16'b00101_001011_00111; 
		4141: oled_colour = 16'b00111_010000_01001; 
		4142: oled_colour = 16'b00011_001010_00111; 
		4143: oled_colour = 16'b00101_001110_01001; 
		4144: oled_colour = 16'b00101_001101_01001; 
		4145: oled_colour = 16'b00100_001001_00111; 
		4146: oled_colour = 16'b00101_001110_01010; 
		4147: oled_colour = 16'b00101_001101_01001; 
		4148: oled_colour = 16'b00100_000111_00101; 
		4149: oled_colour = 16'b00110_001110_01000; 
		4150: oled_colour = 16'b00011_001000_00110; 
		4151: oled_colour = 16'b00101_001100_01000; 
		4152: oled_colour = 16'b00011_000101_00011; 
		4153: oled_colour = 16'b00011_000101_00011; 
		4154: oled_colour = 16'b00011_000101_00011; 
		4155: oled_colour = 16'b00011_000101_00011; 
		4156: oled_colour = 16'b00011_000101_00011; 
		4157: oled_colour = 16'b00010_000100_00011; 
		4158: oled_colour = 16'b00010_000101_00100; 
		4159: oled_colour = 16'b00011_000110_00101; 
		4160: oled_colour = 16'b00011_000111_00101; 
		4161: oled_colour = 16'b00010_000101_00100; 
		4162: oled_colour = 16'b00010_000100_00011; 
		4163: oled_colour = 16'b00100_001000_00100; 
		4164: oled_colour = 16'b00100_000111_00011; 
		4165: oled_colour = 16'b00001_000001_00010; 
		4166: oled_colour = 16'b00010_000101_00100; 
		4167: oled_colour = 16'b01000_010001_01001; 
		4168: oled_colour = 16'b10011_100111_10000; 
		4169: oled_colour = 16'b01101_011100_01100; 
		4170: oled_colour = 16'b10100_101000_10000; 
		4171: oled_colour = 16'b11001_110010_10011; 
		4172: oled_colour = 16'b10001_100100_01111; 
		4173: oled_colour = 16'b01110_011101_01110; 
		4174: oled_colour = 16'b01011_010111_01101; 
		4175: oled_colour = 16'b00110_001110_01001; 
		4176: oled_colour = 16'b01010_010110_01011; 
		4177: oled_colour = 16'b01101_011011_01101; 
		4178: oled_colour = 16'b00110_001110_01001; 
		4179: oled_colour = 16'b01010_010101_01011; 
		4180: oled_colour = 16'b10000_100001_01110; 
		4181: oled_colour = 16'b00111_001111_01001; 
		4182: oled_colour = 16'b01000_010010_01010; 
		4183: oled_colour = 16'b01111_011111_01110; 
		4184: oled_colour = 16'b00111_010000_01010; 
		4185: oled_colour = 16'b00111_010001_01010; 
		4186: oled_colour = 16'b01111_011111_01110; 
		4187: oled_colour = 16'b01000_010010_01010; 
		4188: oled_colour = 16'b00110_001111_01001; 
		4189: oled_colour = 16'b01101_011100_01101; 
		4190: oled_colour = 16'b01001_010011_01011; 
		4191: oled_colour = 16'b00110_001110_01001; 
		4192: oled_colour = 16'b10000_100000_01110; 
		4193: oled_colour = 16'b01011_010111_01011; 
		4194: oled_colour = 16'b00101_001110_01001; 
		4195: oled_colour = 16'b01110_011100_01101; 
		4196: oled_colour = 16'b01011_011000_01100; 
		4197: oled_colour = 16'b00110_001101_01001; 
		4198: oled_colour = 16'b01101_011010_01101; 
		4199: oled_colour = 16'b01101_011011_01100; 
		4200: oled_colour = 16'b00110_001101_01001; 
		4201: oled_colour = 16'b01010_010110_01011; 
		4202: oled_colour = 16'b01101_011011_01101; 
		4203: oled_colour = 16'b00110_001110_01001; 
		4204: oled_colour = 16'b01011_010110_01011; 
		4205: oled_colour = 16'b10001_100010_01111; 
		4206: oled_colour = 16'b00111_001110_01001; 
		4207: oled_colour = 16'b01000_010011_01010; 
		4208: oled_colour = 16'b01111_011111_01110; 
		4209: oled_colour = 16'b00111_010000_01010; 
		4210: oled_colour = 16'b01000_010001_01010; 
		4211: oled_colour = 16'b10000_100000_01110; 
		4212: oled_colour = 16'b01001_010010_01010; 
		4213: oled_colour = 16'b00101_001100_01000; 
		4214: oled_colour = 16'b00101_001110_01000; 
		4215: oled_colour = 16'b00100_001101_01000; 
		4216: oled_colour = 16'b00011_001010_00111; 
		4217: oled_colour = 16'b00100_001100_00111; 
		4218: oled_colour = 16'b00011_001001_00110; 
		4219: oled_colour = 16'b00010_000110_00100; 
		4220: oled_colour = 16'b00011_001000_00101; 
		4221: oled_colour = 16'b00100_001100_01000; 
		4222: oled_colour = 16'b01011_010111_01011; 
		4223: oled_colour = 16'b01101_011011_01100; 
		4224: oled_colour = 16'b00010_000100_00010; 
		4225: oled_colour = 16'b00100_001001_00110; 
		4226: oled_colour = 16'b00101_001100_00111; 
		4227: oled_colour = 16'b00011_000111_00100; 
		4228: oled_colour = 16'b00100_001001_00110; 
		4229: oled_colour = 16'b00101_001011_00111; 
		4230: oled_colour = 16'b00100_001010_00110; 
		4231: oled_colour = 16'b00011_000111_00100; 
		4232: oled_colour = 16'b00100_001001_00110; 
		4233: oled_colour = 16'b00010_000101_00100; 
		4234: oled_colour = 16'b00011_000110_00101; 
		4235: oled_colour = 16'b00100_001010_00111; 
		4236: oled_colour = 16'b00111_010000_01010; 
		4237: oled_colour = 16'b01000_010011_01011; 
		4238: oled_colour = 16'b00010_000100_00100; 
		4239: oled_colour = 16'b00011_001001_00110; 
		4240: oled_colour = 16'b00110_001111_01001; 
		4241: oled_colour = 16'b00100_001001_00110; 
		4242: oled_colour = 16'b00100_001011_00111; 
		4243: oled_colour = 16'b00010_000100_00100; 
		4244: oled_colour = 16'b00110_001101_01000; 
		4245: oled_colour = 16'b01001_010111_01101; 
		4246: oled_colour = 16'b00100_001011_01000; 
		4247: oled_colour = 16'b00011_001000_00110; 
		4248: oled_colour = 16'b00010_000100_00010; 
		4249: oled_colour = 16'b00011_000101_00011; 
		4250: oled_colour = 16'b00011_000101_00011; 
		4251: oled_colour = 16'b00011_000101_00011; 
		4252: oled_colour = 16'b00011_000101_00011; 
		4253: oled_colour = 16'b00011_000101_00010; 
		4254: oled_colour = 16'b00011_000101_00011; 
		4255: oled_colour = 16'b00010_000100_00011; 
		4256: oled_colour = 16'b00010_000101_00011; 
		4257: oled_colour = 16'b00101_001100_00111; 
		4258: oled_colour = 16'b01010_010011_01001; 
		4259: oled_colour = 16'b01110_011100_01011; 
		4260: oled_colour = 16'b01100_011000_01010; 
		4261: oled_colour = 16'b01001_010010_01000; 
		4262: oled_colour = 16'b00101_001010_00101; 
		4263: oled_colour = 16'b00001_000010_00010; 
		4264: oled_colour = 16'b00011_000111_00101; 
		4265: oled_colour = 16'b00100_001011_01000; 
		4266: oled_colour = 16'b01101_011100_01101; 
		4267: oled_colour = 16'b11000_110001_10010; 
		4268: oled_colour = 16'b11101_111000_10100; 
		4269: oled_colour = 16'b11011_110100_10011; 
		4270: oled_colour = 16'b10100_101001_10000; 
		4271: oled_colour = 16'b01100_011011_01101; 
		4272: oled_colour = 16'b01010_010110_01100; 
		4273: oled_colour = 16'b01111_011101_01110; 
		4274: oled_colour = 16'b00110_001110_01001; 
		4275: oled_colour = 16'b01010_010100_01011; 
		4276: oled_colour = 16'b01111_011110_01110; 
		4277: oled_colour = 16'b00111_010000_01010; 
		4278: oled_colour = 16'b01000_010001_01010; 
		4279: oled_colour = 16'b01110_011101_01101; 
		4280: oled_colour = 16'b01000_010001_01010; 
		4281: oled_colour = 16'b01000_010001_01010; 
		4282: oled_colour = 16'b10001_100011_01111; 
		4283: oled_colour = 16'b01001_010011_01011; 
		4284: oled_colour = 16'b00110_001110_01001; 
		4285: oled_colour = 16'b01111_011110_01110; 
		4286: oled_colour = 16'b01001_010100_01011; 
		4287: oled_colour = 16'b00110_001110_01001; 
		4288: oled_colour = 16'b01110_011100_01101; 
		4289: oled_colour = 16'b01011_010110_01011; 
		4290: oled_colour = 16'b00110_001101_01001; 
		4291: oled_colour = 16'b01101_011010_01100; 
		4292: oled_colour = 16'b01100_011000_01100; 
		4293: oled_colour = 16'b00110_001101_01001; 
		4294: oled_colour = 16'b01110_011101_01101; 
		4295: oled_colour = 16'b01111_011110_01110; 
		4296: oled_colour = 16'b00101_001101_01001; 
		4297: oled_colour = 16'b01011_010111_01100; 
		4298: oled_colour = 16'b01111_011110_01110; 
		4299: oled_colour = 16'b00110_001110_01001; 
		4300: oled_colour = 16'b01001_010100_01011; 
		4301: oled_colour = 16'b01111_011110_01110; 
		4302: oled_colour = 16'b00111_001111_01001; 
		4303: oled_colour = 16'b01000_010001_01010; 
		4304: oled_colour = 16'b01111_011110_01101; 
		4305: oled_colour = 16'b00111_010001_01010; 
		4306: oled_colour = 16'b01000_010001_01010; 
		4307: oled_colour = 16'b10010_100011_01111; 
		4308: oled_colour = 16'b01001_010011_01011; 
		4309: oled_colour = 16'b00101_001101_01000; 
		4310: oled_colour = 16'b00110_001111_01001; 
		4311: oled_colour = 16'b00100_001101_01000; 
		4312: oled_colour = 16'b00011_001010_00111; 
		4313: oled_colour = 16'b00011_001010_00111; 
		4314: oled_colour = 16'b00011_001001_00110; 
		4315: oled_colour = 16'b00010_000110_00100; 
		4316: oled_colour = 16'b00011_000110_00100; 
		4317: oled_colour = 16'b00011_001010_00111; 
		4318: oled_colour = 16'b00100_001011_00111; 
		4319: oled_colour = 16'b10011_100110_01111; 
		4320: oled_colour = 16'b00011_000101_00011; 
		4321: oled_colour = 16'b00010_000100_00010; 
		4322: oled_colour = 16'b00011_000110_00100; 
		4323: oled_colour = 16'b00101_001011_00111; 
		4324: oled_colour = 16'b00101_001101_00111; 
		4325: oled_colour = 16'b00101_001011_00111; 
		4326: oled_colour = 16'b00011_000101_00100; 
		4327: oled_colour = 16'b00011_001000_00101; 
		4328: oled_colour = 16'b00100_001010_00110; 
		4329: oled_colour = 16'b00011_001000_00101; 
		4330: oled_colour = 16'b00011_000111_00101; 
		4331: oled_colour = 16'b00100_001010_00111; 
		4332: oled_colour = 16'b00011_001001_00110; 
		4333: oled_colour = 16'b00010_000101_00101; 
		4334: oled_colour = 16'b00110_001101_01000; 
		4335: oled_colour = 16'b00101_001011_00110; 
		4336: oled_colour = 16'b00100_001001_00110; 
		4337: oled_colour = 16'b00111_001110_01000; 
		4338: oled_colour = 16'b00100_001010_00110; 
		4339: oled_colour = 16'b00111_001111_01000; 
		4340: oled_colour = 16'b00100_001000_00101; 
		4341: oled_colour = 16'b00010_000101_00100; 
		4342: oled_colour = 16'b00110_001110_01001; 
		4343: oled_colour = 16'b01001_010100_01010; 
		4344: oled_colour = 16'b00011_000111_00101; 
		4345: oled_colour = 16'b00010_000011_00010; 
		4346: oled_colour = 16'b00010_000100_00010; 
		4347: oled_colour = 16'b00011_000101_00011; 
		4348: oled_colour = 16'b00011_000101_00011; 
		4349: oled_colour = 16'b00011_000101_00011; 
		4350: oled_colour = 16'b00010_000100_00010; 
		4351: oled_colour = 16'b00011_000110_00100; 
		4352: oled_colour = 16'b00111_001110_01000; 
		4353: oled_colour = 16'b01001_010011_01001; 
		4354: oled_colour = 16'b00101_001100_00111; 
		4355: oled_colour = 16'b01000_010010_01010; 
		4356: oled_colour = 16'b00111_010001_01001; 
		4357: oled_colour = 16'b00110_001101_00111; 
		4358: oled_colour = 16'b01001_010011_01001; 
		4359: oled_colour = 16'b00110_001101_00111; 
		4360: oled_colour = 16'b00011_000101_00011; 
		4361: oled_colour = 16'b00010_000100_00011; 
		4362: oled_colour = 16'b00011_000111_00101; 
		4363: oled_colour = 16'b00111_010001_01010; 
		4364: oled_colour = 16'b01111_011111_01110; 
		4365: oled_colour = 16'b10110_101101_10001; 
		4366: oled_colour = 16'b11110_111001_10100; 
		4367: oled_colour = 16'b10000_100000_01101; 
		4368: oled_colour = 16'b01100_011011_01100; 
		4369: oled_colour = 16'b01111_100000_01110; 
		4370: oled_colour = 16'b00110_001111_01010; 
		4371: oled_colour = 16'b01000_010011_01011; 
		4372: oled_colour = 16'b01111_011111_01110; 
		4373: oled_colour = 16'b00110_001110_01001; 
		4374: oled_colour = 16'b01000_010001_01010; 
		4375: oled_colour = 16'b01111_011111_01110; 
		4376: oled_colour = 16'b00111_010000_01010; 
		4377: oled_colour = 16'b00111_010000_01010; 
		4378: oled_colour = 16'b10000_100000_01110; 
		4379: oled_colour = 16'b01001_010010_01010; 
		4380: oled_colour = 16'b00110_001110_01001; 
		4381: oled_colour = 16'b01111_011111_01110; 
		4382: oled_colour = 16'b01001_010011_01010; 
		4383: oled_colour = 16'b00110_001110_01001; 
		4384: oled_colour = 16'b01110_011101_01101; 
		4385: oled_colour = 16'b01010_010110_01011; 
		4386: oled_colour = 16'b00101_001100_01000; 
		4387: oled_colour = 16'b01110_011101_01101; 
		4388: oled_colour = 16'b01100_011001_01100; 
		4389: oled_colour = 16'b00101_001100_01000; 
		4390: oled_colour = 16'b01101_011011_01101; 
		4391: oled_colour = 16'b01110_011100_01101; 
		4392: oled_colour = 16'b00101_001100_01000; 
		4393: oled_colour = 16'b01011_011000_01100; 
		4394: oled_colour = 16'b01111_011110_01101; 
		4395: oled_colour = 16'b00110_001101_01001; 
		4396: oled_colour = 16'b01001_010100_01011; 
		4397: oled_colour = 16'b01111_011111_01110; 
		4398: oled_colour = 16'b00110_001110_01001; 
		4399: oled_colour = 16'b01000_010010_01010; 
		4400: oled_colour = 16'b10000_100000_01110; 
		4401: oled_colour = 16'b00111_010001_01010; 
		4402: oled_colour = 16'b00111_010000_01001; 
		4403: oled_colour = 16'b10000_100001_01110; 
		4404: oled_colour = 16'b01001_010010_01010; 
		4405: oled_colour = 16'b00101_001101_01000; 
		4406: oled_colour = 16'b00110_001111_01001; 
		4407: oled_colour = 16'b00100_001101_01000; 
		4408: oled_colour = 16'b00011_001010_00111; 
		4409: oled_colour = 16'b00100_001010_00111; 
		4410: oled_colour = 16'b00011_001000_00101; 
		4411: oled_colour = 16'b00010_000101_00011; 
		4412: oled_colour = 16'b00011_000110_00100; 
		4413: oled_colour = 16'b00011_001010_00111; 
		4414: oled_colour = 16'b00011_001001_00111; 
		4415: oled_colour = 16'b01111_011110_01101; 
		4416: oled_colour = 16'b00011_000111_00101; 
		4417: oled_colour = 16'b00011_000100_00011; 
		4418: oled_colour = 16'b00010_000100_00011; 
		4419: oled_colour = 16'b00010_000100_00010; 
		4420: oled_colour = 16'b00011_000111_00100; 
		4421: oled_colour = 16'b00101_001011_00111; 
		4422: oled_colour = 16'b00110_001101_00111; 
		4423: oled_colour = 16'b00110_001110_01000; 
		4424: oled_colour = 16'b00101_001100_00110; 
		4425: oled_colour = 16'b00110_001101_00110; 
		4426: oled_colour = 16'b00110_001101_01000; 
		4427: oled_colour = 16'b00101_001101_01000; 
		4428: oled_colour = 16'b00101_001011_00111; 
		4429: oled_colour = 16'b00011_000101_00100; 
		4430: oled_colour = 16'b00111_010001_01010; 
		4431: oled_colour = 16'b00110_001111_01001; 
		4432: oled_colour = 16'b00011_000111_00101; 
		4433: oled_colour = 16'b01000_010001_01001; 
		4434: oled_colour = 16'b00100_001001_00110; 
		4435: oled_colour = 16'b00111_010010_01011; 
		4436: oled_colour = 16'b00100_001001_00110; 
		4437: oled_colour = 16'b00011_001000_00101; 
		4438: oled_colour = 16'b00110_001101_01000; 
		4439: oled_colour = 16'b10010_100101_10000; 
		4440: oled_colour = 16'b10000_100010_01111; 
		4441: oled_colour = 16'b01000_010010_01001; 
		4442: oled_colour = 16'b00100_001001_00101; 
		4443: oled_colour = 16'b00010_000101_00011; 
		4444: oled_colour = 16'b00010_000100_00010; 
		4445: oled_colour = 16'b00011_000100_00010; 
		4446: oled_colour = 16'b00011_000101_00011; 
		4447: oled_colour = 16'b00101_001011_00111; 
		4448: oled_colour = 16'b00011_001000_00110; 
		4449: oled_colour = 16'b01001_010101_01011; 
		4450: oled_colour = 16'b01000_010011_01011; 
		4451: oled_colour = 16'b00101_001110_01001; 
		4452: oled_colour = 16'b00101_001110_01001; 
		4453: oled_colour = 16'b01000_010011_01011; 
		4454: oled_colour = 16'b00111_010001_01010; 
		4455: oled_colour = 16'b00011_001001_00110; 
		4456: oled_colour = 16'b00100_001010_00111; 
		4457: oled_colour = 16'b00011_000101_00011; 
		4458: oled_colour = 16'b00010_000100_00010; 
		4459: oled_colour = 16'b00010_000100_00011; 
		4460: oled_colour = 16'b00011_000110_00101; 
		4461: oled_colour = 16'b00111_010000_01001; 
		4462: oled_colour = 16'b01110_011110_01110; 
		4463: oled_colour = 16'b01000_010010_01001; 
		4464: oled_colour = 16'b10101_101001_10001; 
		4465: oled_colour = 16'b11010_110011_10011; 
		4466: oled_colour = 16'b10011_100111_10000; 
		4467: oled_colour = 16'b01110_011101_01110; 
		4468: oled_colour = 16'b01100_011011_01101; 
		4469: oled_colour = 16'b01000_010010_01011; 
		4470: oled_colour = 16'b01000_010011_01011; 
		4471: oled_colour = 16'b10001_100001_01110; 
		4472: oled_colour = 16'b01000_010000_01010; 
		4473: oled_colour = 16'b00111_010000_01010; 
		4474: oled_colour = 16'b01111_011110_01110; 
		4475: oled_colour = 16'b01000_010010_01010; 
		4476: oled_colour = 16'b00111_010000_01010; 
		4477: oled_colour = 16'b10001_100010_01111; 
		4478: oled_colour = 16'b01001_010100_01010; 
		4479: oled_colour = 16'b00110_001110_01001; 
		4480: oled_colour = 16'b01110_011101_01101; 
		4481: oled_colour = 16'b01010_010111_01011; 
		4482: oled_colour = 16'b00101_001100_01001; 
		4483: oled_colour = 16'b01111_011111_01110; 
		4484: oled_colour = 16'b01101_011010_01100; 
		4485: oled_colour = 16'b00101_001100_01001; 
		4486: oled_colour = 16'b01100_011001_01100; 
		4487: oled_colour = 16'b01101_011011_01101; 
		4488: oled_colour = 16'b00101_001100_01001; 
		4489: oled_colour = 16'b01101_011010_01101; 
		4490: oled_colour = 16'b10000_011111_01110; 
		4491: oled_colour = 16'b00110_001101_01001; 
		4492: oled_colour = 16'b01001_010100_01011; 
		4493: oled_colour = 16'b01111_011111_01110; 
		4494: oled_colour = 16'b00110_001111_01001; 
		4495: oled_colour = 16'b01000_010011_01010; 
		4496: oled_colour = 16'b10001_100010_01110; 
		4497: oled_colour = 16'b00111_010000_01010; 
		4498: oled_colour = 16'b00111_010000_01010; 
		4499: oled_colour = 16'b01111_011111_01101; 
		4500: oled_colour = 16'b01000_010011_01010; 
		4501: oled_colour = 16'b00110_001111_01001; 
		4502: oled_colour = 16'b01000_010001_01010; 
		4503: oled_colour = 16'b00101_001101_01000; 
		4504: oled_colour = 16'b00011_001010_00111; 
		4505: oled_colour = 16'b00100_001010_00111; 
		4506: oled_colour = 16'b00011_001000_00110; 
		4507: oled_colour = 16'b00010_000110_00011; 
		4508: oled_colour = 16'b00011_000110_00100; 
		4509: oled_colour = 16'b00011_001010_00111; 
		4510: oled_colour = 16'b00010_001001_00111; 
		4511: oled_colour = 16'b00101_001101_01000; 
		4512: oled_colour = 16'b00011_001001_00111; 
		4513: oled_colour = 16'b00010_000101_00011; 
		4514: oled_colour = 16'b00011_000100_00011; 
		4515: oled_colour = 16'b00011_000101_00011; 
		4516: oled_colour = 16'b00010_000100_00010; 
		4517: oled_colour = 16'b00010_000100_00010; 
		4518: oled_colour = 16'b00011_000101_00011; 
		4519: oled_colour = 16'b00011_000110_00100; 
		4520: oled_colour = 16'b00100_001001_00101; 
		4521: oled_colour = 16'b00100_001000_00101; 
		4522: oled_colour = 16'b00100_001000_00101; 
		4523: oled_colour = 16'b00010_000100_00010; 
		4524: oled_colour = 16'b00011_000111_00100; 
		4525: oled_colour = 16'b00101_001011_00111; 
		4526: oled_colour = 16'b00011_001000_00110; 
		4527: oled_colour = 16'b00010_000101_00011; 
		4528: oled_colour = 16'b00100_001001_00110; 
		4529: oled_colour = 16'b00110_001110_01001; 
		4530: oled_colour = 16'b00010_000100_00011; 
		4531: oled_colour = 16'b00010_000101_00100; 
		4532: oled_colour = 16'b00100_001010_00110; 
		4533: oled_colour = 16'b00100_001010_00111; 
		4534: oled_colour = 16'b00010_000110_00101; 
		4535: oled_colour = 16'b00111_001110_01001; 
		4536: oled_colour = 16'b10101_101010_10001; 
		4537: oled_colour = 16'b10101_101011_10000; 
		4538: oled_colour = 16'b01110_011110_01110; 
		4539: oled_colour = 16'b00111_010001_01010; 
		4540: oled_colour = 16'b00100_001001_00110; 
		4541: oled_colour = 16'b00010_000011_00011; 
		4542: oled_colour = 16'b00100_001001_00110; 
		4543: oled_colour = 16'b00101_001101_01000; 
		4544: oled_colour = 16'b00100_001100_01000; 
		4545: oled_colour = 16'b00100_001000_00110; 
		4546: oled_colour = 16'b00100_001010_00111; 
		4547: oled_colour = 16'b00100_001001_00101; 
		4548: oled_colour = 16'b00011_000110_00101; 
		4549: oled_colour = 16'b00100_001001_00111; 
		4550: oled_colour = 16'b00011_000111_00110; 
		4551: oled_colour = 16'b00101_001110_01001; 
		4552: oled_colour = 16'b00110_001110_01000; 
		4553: oled_colour = 16'b00100_001010_00111; 
		4554: oled_colour = 16'b00011_000110_00100; 
		4555: oled_colour = 16'b00011_000101_00011; 
		4556: oled_colour = 16'b00010_000100_00010; 
		4557: oled_colour = 16'b00010_000100_00011; 
		4558: oled_colour = 16'b00010_000101_00100; 
		4559: oled_colour = 16'b00011_001000_00111; 
		4560: oled_colour = 16'b01001_010110_01100; 
		4561: oled_colour = 16'b10100_101001_10001; 
		4562: oled_colour = 16'b11100_110101_10011; 
		4563: oled_colour = 16'b11011_110100_10011; 
		4564: oled_colour = 16'b10110_101100_10001; 
		4565: oled_colour = 16'b01011_011001_01100; 
		4566: oled_colour = 16'b00101_001101_01001; 
		4567: oled_colour = 16'b01101_011011_01101; 
		4568: oled_colour = 16'b01000_010001_01010; 
		4569: oled_colour = 16'b00111_010000_01010; 
		4570: oled_colour = 16'b01110_011101_01101; 
		4571: oled_colour = 16'b01001_010011_01010; 
		4572: oled_colour = 16'b00110_001110_01001; 
		4573: oled_colour = 16'b01111_011110_01110; 
		4574: oled_colour = 16'b01001_010011_01011; 
		4575: oled_colour = 16'b00110_001110_01001; 
		4576: oled_colour = 16'b01111_011110_01101; 
		4577: oled_colour = 16'b01011_010111_01011; 
		4578: oled_colour = 16'b00110_001101_01001; 
		4579: oled_colour = 16'b01100_011010_01100; 
		4580: oled_colour = 16'b01011_010111_01011; 
		4581: oled_colour = 16'b00110_001101_01001; 
		4582: oled_colour = 16'b01011_011000_01100; 
		4583: oled_colour = 16'b01101_011010_01101; 
		4584: oled_colour = 16'b00110_001101_01001; 
		4585: oled_colour = 16'b01011_010111_01100; 
		4586: oled_colour = 16'b01111_011101_01110; 
		4587: oled_colour = 16'b00110_001110_01001; 
		4588: oled_colour = 16'b01001_010101_01011; 
		4589: oled_colour = 16'b10000_100000_01110; 
		4590: oled_colour = 16'b00111_010000_01010; 
		4591: oled_colour = 16'b01000_010001_01010; 
		4592: oled_colour = 16'b01110_011100_01101; 
		4593: oled_colour = 16'b01000_010001_01010; 
		4594: oled_colour = 16'b00111_001111_01010; 
		4595: oled_colour = 16'b01111_011110_01101; 
		4596: oled_colour = 16'b01001_010011_01010; 
		4597: oled_colour = 16'b00110_001111_01001; 
		4598: oled_colour = 16'b00111_010000_01010; 
		4599: oled_colour = 16'b00100_001101_01000; 
		4600: oled_colour = 16'b00011_001010_00111; 
		4601: oled_colour = 16'b00100_001011_00111; 
		4602: oled_colour = 16'b00011_001001_00110; 
		4603: oled_colour = 16'b00010_000110_00100; 
		4604: oled_colour = 16'b00011_000110_00100; 
		4605: oled_colour = 16'b00011_001001_00110; 
		4606: oled_colour = 16'b00011_001001_00110; 
		4607: oled_colour = 16'b00010_000101_00100; 
		4608: oled_colour = 16'b00101_001110_01001; 
		4609: oled_colour = 16'b00100_001010_00111; 
		4610: oled_colour = 16'b00010_000100_00011; 
		4611: oled_colour = 16'b00011_000100_00010; 
		4612: oled_colour = 16'b00011_000101_00011; 
		4613: oled_colour = 16'b00011_000101_00011; 
		4614: oled_colour = 16'b00011_000101_00011; 
		4615: oled_colour = 16'b00010_000100_00010; 
		4616: oled_colour = 16'b00010_000100_00010; 
		4617: oled_colour = 16'b00010_000100_00010; 
		4618: oled_colour = 16'b00010_000100_00010; 
		4619: oled_colour = 16'b00011_000101_00010; 
		4620: oled_colour = 16'b00010_000100_00010; 
		4621: oled_colour = 16'b00011_000101_00011; 
		4622: oled_colour = 16'b00100_001001_00110; 
		4623: oled_colour = 16'b00101_001100_00111; 
		4624: oled_colour = 16'b00110_001110_00111; 
		4625: oled_colour = 16'b00111_001110_01000; 
		4626: oled_colour = 16'b00110_001101_00111; 
		4627: oled_colour = 16'b00100_001011_00111; 
		4628: oled_colour = 16'b00011_000111_00101; 
		4629: oled_colour = 16'b00011_000100_00011; 
		4630: oled_colour = 16'b01010_010111_01100; 
		4631: oled_colour = 16'b00110_010001_01010; 
		4632: oled_colour = 16'b00100_001011_01000; 
		4633: oled_colour = 16'b10001_100010_01111; 
		4634: oled_colour = 16'b10110_101100_10001; 
		4635: oled_colour = 16'b10100_101001_10000; 
		4636: oled_colour = 16'b10001_100100_01111; 
		4637: oled_colour = 16'b01110_011101_01101; 
		4638: oled_colour = 16'b00100_001011_00111; 
		4639: oled_colour = 16'b00101_001101_01000; 
		4640: oled_colour = 16'b00100_001100_01000; 
		4641: oled_colour = 16'b00100_001001_00110; 
		4642: oled_colour = 16'b01001_010101_01011; 
		4643: oled_colour = 16'b01001_010100_01011; 
		4644: oled_colour = 16'b00101_001100_01000; 
		4645: oled_colour = 16'b00100_001011_00111; 
		4646: oled_colour = 16'b00100_001011_00111; 
		4647: oled_colour = 16'b01000_010010_01011; 
		4648: oled_colour = 16'b00110_001110_01001; 
		4649: oled_colour = 16'b00100_001001_00111; 
		4650: oled_colour = 16'b00011_000111_00101; 
		4651: oled_colour = 16'b00011_000110_00101; 
		4652: oled_colour = 16'b00011_000110_00100; 
		4653: oled_colour = 16'b00011_000101_00011; 
		4654: oled_colour = 16'b00011_000100_00010; 
		4655: oled_colour = 16'b00010_000100_00011; 
		4656: oled_colour = 16'b00010_000110_00101; 
		4657: oled_colour = 16'b00101_001100_01000; 
		4658: oled_colour = 16'b01011_011000_01101; 
		4659: oled_colour = 16'b10101_101011_10001; 
		4660: oled_colour = 16'b11100_110110_10011; 
		4661: oled_colour = 16'b01110_011100_01100; 
		4662: oled_colour = 16'b10011_100111_10000; 
		4663: oled_colour = 16'b10000_100001_01111; 
		4664: oled_colour = 16'b01000_010010_01011; 
		4665: oled_colour = 16'b00111_010000_01010; 
		4666: oled_colour = 16'b01111_011111_01110; 
		4667: oled_colour = 16'b01000_010010_01010; 
		4668: oled_colour = 16'b00110_001111_01001; 
		4669: oled_colour = 16'b01110_011100_01101; 
		4670: oled_colour = 16'b01001_010100_01011; 
		4671: oled_colour = 16'b00110_001111_01010; 
		4672: oled_colour = 16'b01101_011011_01101; 
		4673: oled_colour = 16'b01010_010101_01011; 
		4674: oled_colour = 16'b00101_001101_01001; 
		4675: oled_colour = 16'b01101_011100_01101; 
		4676: oled_colour = 16'b01100_011001_01100; 
		4677: oled_colour = 16'b00110_001110_01001; 
		4678: oled_colour = 16'b01101_011011_01101; 
		4679: oled_colour = 16'b01101_011011_01101; 
		4680: oled_colour = 16'b00110_001101_01001; 
		4681: oled_colour = 16'b01011_010110_01011; 
		4682: oled_colour = 16'b01101_011100_01101; 
		4683: oled_colour = 16'b00110_001111_01001; 
		4684: oled_colour = 16'b01001_010100_01011; 
		4685: oled_colour = 16'b01101_011100_01101; 
		4686: oled_colour = 16'b00110_001111_01001; 
		4687: oled_colour = 16'b01000_010001_01010; 
		4688: oled_colour = 16'b01111_011111_01110; 
		4689: oled_colour = 16'b01000_010010_01010; 
		4690: oled_colour = 16'b01000_010001_01010; 
		4691: oled_colour = 16'b10000_100000_01110; 
		4692: oled_colour = 16'b01000_010010_01010; 
		4693: oled_colour = 16'b00111_010000_01001; 
		4694: oled_colour = 16'b01000_010010_01010; 
		4695: oled_colour = 16'b00100_001100_01000; 
		4696: oled_colour = 16'b00100_001011_00111; 
		4697: oled_colour = 16'b00011_001001_00111; 
		4698: oled_colour = 16'b00011_001000_00110; 
		4699: oled_colour = 16'b00010_000110_00100; 
		4700: oled_colour = 16'b00011_000111_00100; 
		4701: oled_colour = 16'b00010_000110_00100; 
		4702: oled_colour = 16'b00010_000101_00011; 
		4703: oled_colour = 16'b00111_001110_01000; 
		4704: oled_colour = 16'b00101_001010_00110; 
		4705: oled_colour = 16'b00110_001111_01001; 
		4706: oled_colour = 16'b00100_001001_00111; 
		4707: oled_colour = 16'b00011_000101_00011; 
		4708: oled_colour = 16'b00010_000100_00010; 
		4709: oled_colour = 16'b00011_000101_00011; 
		4710: oled_colour = 16'b00011_000101_00011; 
		4711: oled_colour = 16'b00011_000101_00011; 
		4712: oled_colour = 16'b00011_000101_00011; 
		4713: oled_colour = 16'b00011_000101_00011; 
		4714: oled_colour = 16'b00011_000101_00011; 
		4715: oled_colour = 16'b00011_000101_00011; 
		4716: oled_colour = 16'b00011_000101_00011; 
		4717: oled_colour = 16'b00011_000101_00010; 
		4718: oled_colour = 16'b00010_000100_00010; 
		4719: oled_colour = 16'b00011_000101_00011; 
		4720: oled_colour = 16'b00100_001010_00110; 
		4721: oled_colour = 16'b00110_001101_00111; 
		4722: oled_colour = 16'b00011_000111_00101; 
		4723: oled_colour = 16'b00010_000101_00011; 
		4724: oled_colour = 16'b00011_000100_00011; 
		4725: oled_colour = 16'b00011_000101_00011; 
		4726: oled_colour = 16'b01100_011010_01101; 
		4727: oled_colour = 16'b10100_101010_10001; 
		4728: oled_colour = 16'b01100_011001_01100; 
		4729: oled_colour = 16'b00100_001011_01000; 
		4730: oled_colour = 16'b00101_001101_01000; 
		4731: oled_colour = 16'b01010_010111_01011; 
		4732: oled_colour = 16'b01111_011111_01101; 
		4733: oled_colour = 16'b01111_011111_01110; 
		4734: oled_colour = 16'b00011_001000_00110; 
		4735: oled_colour = 16'b00011_000110_00101; 
		4736: oled_colour = 16'b00011_000110_00100; 
		4737: oled_colour = 16'b00101_001100_00111; 
		4738: oled_colour = 16'b00101_001101_01000; 
		4739: oled_colour = 16'b00101_001110_01001; 
		4740: oled_colour = 16'b00100_001011_01000; 
		4741: oled_colour = 16'b00011_001000_00110; 
		4742: oled_colour = 16'b00101_001100_01000; 
		4743: oled_colour = 16'b00011_001000_00111; 
		4744: oled_colour = 16'b00011_001000_00110; 
		4745: oled_colour = 16'b00011_001001_00110; 
		4746: oled_colour = 16'b00011_000111_00101; 
		4747: oled_colour = 16'b00010_000100_00011; 
		4748: oled_colour = 16'b00011_000110_00101; 
		4749: oled_colour = 16'b00011_000110_00101; 
		4750: oled_colour = 16'b00011_000111_00100; 
		4751: oled_colour = 16'b00011_000110_00011; 
		4752: oled_colour = 16'b00011_000101_00010; 
		4753: oled_colour = 16'b00010_000100_00011; 
		4754: oled_colour = 16'b00010_000110_00101; 
		4755: oled_colour = 16'b00110_001110_01001; 
		4756: oled_colour = 16'b01010_010110_01011; 
		4757: oled_colour = 16'b01001_010100_01010; 
		4758: oled_colour = 16'b11000_110000_10010; 
		4759: oled_colour = 16'b11010_110100_10011; 
		4760: oled_colour = 16'b10111_101100_10001; 
		4761: oled_colour = 16'b10001_100011_01111; 
		4762: oled_colour = 16'b01110_011101_01110; 
		4763: oled_colour = 16'b01001_010101_01011; 
		4764: oled_colour = 16'b00111_010001_01011; 
		4765: oled_colour = 16'b01111_011110_01110; 
		4766: oled_colour = 16'b01010_010100_01011; 
		4767: oled_colour = 16'b00111_001111_01010; 
		4768: oled_colour = 16'b01100_011001_01100; 
		4769: oled_colour = 16'b01010_010101_01011; 
		4770: oled_colour = 16'b00110_001101_01001; 
		4771: oled_colour = 16'b01110_011110_01101; 
		4772: oled_colour = 16'b01101_011011_01100; 
		4773: oled_colour = 16'b00110_001110_01001; 
		4774: oled_colour = 16'b01011_011000_01100; 
		4775: oled_colour = 16'b01100_011010_01100; 
		4776: oled_colour = 16'b00110_001110_01001; 
		4777: oled_colour = 16'b01011_010111_01100; 
		4778: oled_colour = 16'b01110_011101_01110; 
		4779: oled_colour = 16'b00111_001111_01010; 
		4780: oled_colour = 16'b01001_010011_01011; 
		4781: oled_colour = 16'b01101_011011_01101; 
		4782: oled_colour = 16'b00111_010000_01001; 
		4783: oled_colour = 16'b01000_010010_01010; 
		4784: oled_colour = 16'b10001_100010_01110; 
		4785: oled_colour = 16'b01001_010010_01010; 
		4786: oled_colour = 16'b01000_010001_01010; 
		4787: oled_colour = 16'b01110_011100_01101; 
		4788: oled_colour = 16'b01001_010011_01010; 
		4789: oled_colour = 16'b00111_010000_01001; 
		4790: oled_colour = 16'b01100_011001_01100; 
		4791: oled_colour = 16'b00101_001110_01000; 
		4792: oled_colour = 16'b00100_001011_00111; 
		4793: oled_colour = 16'b00011_001001_00110; 
		4794: oled_colour = 16'b00011_001000_00110; 
		4795: oled_colour = 16'b00010_000101_00011; 
		4796: oled_colour = 16'b00010_000101_00100; 
		4797: oled_colour = 16'b00100_001001_00110; 
		4798: oled_colour = 16'b00110_001100_00111; 
		4799: oled_colour = 16'b01100_011010_01101; 
		4800: oled_colour = 16'b00010_000011_00010; 
		4801: oled_colour = 16'b00010_000100_00011; 
		4802: oled_colour = 16'b00011_001000_00101; 
		4803: oled_colour = 16'b00101_001100_01000; 
		4804: oled_colour = 16'b00011_001000_00101; 
		4805: oled_colour = 16'b00010_000100_00010; 
		4806: oled_colour = 16'b00010_000100_00011; 
		4807: oled_colour = 16'b00010_000100_00011; 
		4808: oled_colour = 16'b00010_000100_00011; 
		4809: oled_colour = 16'b00010_000100_00011; 
		4810: oled_colour = 16'b00010_000100_00011; 
		4811: oled_colour = 16'b00010_000100_00011; 
		4812: oled_colour = 16'b00010_000100_00011; 
		4813: oled_colour = 16'b00010_000100_00011; 
		4814: oled_colour = 16'b00010_000100_00011; 
		4815: oled_colour = 16'b00010_000100_00010; 
		4816: oled_colour = 16'b00001_000011_00010; 
		4817: oled_colour = 16'b00001_000010_00010; 
		4818: oled_colour = 16'b00010_000101_00011; 
		4819: oled_colour = 16'b00010_000110_00101; 
		4820: oled_colour = 16'b00011_000101_00101; 
		4821: oled_colour = 16'b00010_000100_00011; 
		4822: oled_colour = 16'b00010_000110_00100; 
		4823: oled_colour = 16'b01111_011110_01101; 
		4824: oled_colour = 16'b10111_101111_10010; 
		4825: oled_colour = 16'b10011_100111_10000; 
		4826: oled_colour = 16'b01100_011011_01101; 
		4827: oled_colour = 16'b00111_010001_01010; 
		4828: oled_colour = 16'b00100_001011_01000; 
		4829: oled_colour = 16'b00011_001001_00111; 
		4830: oled_colour = 16'b00011_000111_00110; 
		4831: oled_colour = 16'b00011_000110_00110; 
		4832: oled_colour = 16'b00010_000101_00100; 
		4833: oled_colour = 16'b00010_000101_00101; 
		4834: oled_colour = 16'b00011_000111_00110; 
		4835: oled_colour = 16'b00011_001000_00110; 
		4836: oled_colour = 16'b00011_001000_00110; 
		4837: oled_colour = 16'b00100_001001_00111; 
		4838: oled_colour = 16'b00010_000111_00110; 
		4839: oled_colour = 16'b00010_000111_00110; 
		4840: oled_colour = 16'b00100_001011_01000; 
		4841: oled_colour = 16'b00011_000111_00110; 
		4842: oled_colour = 16'b00011_000111_00101; 
		4843: oled_colour = 16'b00010_000011_00010; 
		4844: oled_colour = 16'b00010_000100_00011; 
		4845: oled_colour = 16'b00010_000100_00011; 
		4846: oled_colour = 16'b00010_000101_00101; 
		4847: oled_colour = 16'b00011_000110_00101; 
		4848: oled_colour = 16'b00011_000110_00100; 
		4849: oled_colour = 16'b00010_000101_00011; 
		4850: oled_colour = 16'b00010_000100_00010; 
		4851: oled_colour = 16'b00001_000011_00010; 
		4852: oled_colour = 16'b00001_000011_00011; 
		4853: oled_colour = 16'b00010_000100_00100; 
		4854: oled_colour = 16'b00100_001011_01000; 
		4855: oled_colour = 16'b01111_011111_01110; 
		4856: oled_colour = 16'b11001_110010_10011; 
		4857: oled_colour = 16'b11101_111000_10100; 
		4858: oled_colour = 16'b11010_110011_10011; 
		4859: oled_colour = 16'b10101_101010_10001; 
		4860: oled_colour = 16'b01100_011010_01101; 
		4861: oled_colour = 16'b01101_011011_01101; 
		4862: oled_colour = 16'b01001_010100_01011; 
		4863: oled_colour = 16'b00101_001110_01010; 
		4864: oled_colour = 16'b01110_011110_01110; 
		4865: oled_colour = 16'b01011_010111_01100; 
		4866: oled_colour = 16'b00110_001110_01001; 
		4867: oled_colour = 16'b01101_011100_01101; 
		4868: oled_colour = 16'b01100_011001_01100; 
		4869: oled_colour = 16'b00110_001111_01010; 
		4870: oled_colour = 16'b01011_011000_01100; 
		4871: oled_colour = 16'b01100_011001_01100; 
		4872: oled_colour = 16'b00110_001110_01010; 
		4873: oled_colour = 16'b01011_011000_01100; 
		4874: oled_colour = 16'b01110_011101_01110; 
		4875: oled_colour = 16'b00110_001101_01001; 
		4876: oled_colour = 16'b01001_010101_01011; 
		4877: oled_colour = 16'b01111_100000_01110; 
		4878: oled_colour = 16'b00111_010000_01010; 
		4879: oled_colour = 16'b01000_010010_01010; 
		4880: oled_colour = 16'b01111_011111_01110; 
		4881: oled_colour = 16'b01000_010010_01010; 
		4882: oled_colour = 16'b00111_010000_01010; 
		4883: oled_colour = 16'b01101_011100_01101; 
		4884: oled_colour = 16'b01000_010011_01011; 
		4885: oled_colour = 16'b00110_001111_01010; 
		4886: oled_colour = 16'b01110_011101_01110; 
		4887: oled_colour = 16'b00110_010000_01001; 
		4888: oled_colour = 16'b00011_001001_00111; 
		4889: oled_colour = 16'b00100_001010_00111; 
		4890: oled_colour = 16'b00100_001011_00111; 
		4891: oled_colour = 16'b00110_001110_01000; 
		4892: oled_colour = 16'b01011_011000_01101; 
		4893: oled_colour = 16'b10100_101001_10001; 
		4894: oled_colour = 16'b10111_101101_10010; 
		4895: oled_colour = 16'b01001_010100_01010; 
		4896: oled_colour = 16'b00101_000111_00010; 
		4897: oled_colour = 16'b00101_000111_00010; 
		4898: oled_colour = 16'b00101_000111_00010; 
		4899: oled_colour = 16'b00110_001000_00011; 
		4900: oled_colour = 16'b00111_001100_00101; 
		4901: oled_colour = 16'b00111_001100_00101; 
		4902: oled_colour = 16'b00110_001000_00011; 
		4903: oled_colour = 16'b00110_001000_00010; 
		4904: oled_colour = 16'b00101_000111_00010; 
		4905: oled_colour = 16'b00101_001000_00010; 
		4906: oled_colour = 16'b00101_000111_00010; 
		4907: oled_colour = 16'b00101_001000_00011; 
		4908: oled_colour = 16'b00101_000111_00010; 
		4909: oled_colour = 16'b00110_001000_00010; 
		4910: oled_colour = 16'b00101_000111_00010; 
		4911: oled_colour = 16'b00101_000111_00010; 
		4912: oled_colour = 16'b00110_001010_00011; 
		4913: oled_colour = 16'b00110_001001_00010; 
		4914: oled_colour = 16'b00110_001001_00011; 
		4915: oled_colour = 16'b00110_001001_00011; 
		4916: oled_colour = 16'b00101_001000_00010; 
		4917: oled_colour = 16'b00110_001001_00011; 
		4918: oled_colour = 16'b00110_001000_00010; 
		4919: oled_colour = 16'b00100_000110_00010; 
		4920: oled_colour = 16'b01001_010001_00111; 
		4921: oled_colour = 16'b10001_011111_01011; 
		4922: oled_colour = 16'b10110_101000_01110; 
		4923: oled_colour = 16'b10100_100110_01101; 
		4924: oled_colour = 16'b10010_100010_01100; 
		4925: oled_colour = 16'b01010_010011_00111; 
		4926: oled_colour = 16'b00100_000110_00010; 
		4927: oled_colour = 16'b00110_001000_00011; 
		4928: oled_colour = 16'b00110_001000_00010; 
		4929: oled_colour = 16'b00110_001000_00010; 
		4930: oled_colour = 16'b00110_001010_00100; 
		4931: oled_colour = 16'b00110_001000_00011; 
		4932: oled_colour = 16'b00110_001000_00011; 
		4933: oled_colour = 16'b00110_001010_00100; 
		4934: oled_colour = 16'b00110_001000_00011; 
		4935: oled_colour = 16'b00101_001000_00010; 
		4936: oled_colour = 16'b00101_001000_00010; 
		4937: oled_colour = 16'b00101_001000_00010; 
		4938: oled_colour = 16'b00101_001000_00011; 
		4939: oled_colour = 16'b00101_000111_00010; 
		4940: oled_colour = 16'b00110_001000_00010; 
		4941: oled_colour = 16'b00110_001000_00010; 
		4942: oled_colour = 16'b00110_001000_00010; 
		4943: oled_colour = 16'b00101_000111_00010; 
		4944: oled_colour = 16'b00101_000111_00011; 
		4945: oled_colour = 16'b00110_001001_00100; 
		4946: oled_colour = 16'b00110_001010_00100; 
		4947: oled_colour = 16'b00110_001001_00010; 
		4948: oled_colour = 16'b00110_001000_00010; 
		4949: oled_colour = 16'b00101_000111_00010; 
		4950: oled_colour = 16'b00101_000111_00010; 
		4951: oled_colour = 16'b00101_001000_00100; 
		4952: oled_colour = 16'b01010_010001_00111; 
		4953: oled_colour = 16'b10011_100010_01100; 
		4954: oled_colour = 16'b11010_110001_10000; 
		4955: oled_colour = 16'b11100_110011_10001; 
		4956: oled_colour = 16'b10001_011111_01011; 
		4957: oled_colour = 16'b10000_011111_01100; 
		4958: oled_colour = 16'b01111_011100_01011; 
		4959: oled_colour = 16'b01011_010100_01001; 
		4960: oled_colour = 16'b01101_011001_01010; 
		4961: oled_colour = 16'b01110_011001_01010; 
		4962: oled_colour = 16'b01011_010101_01000; 
		4963: oled_colour = 16'b10000_011101_01011; 
		4964: oled_colour = 16'b01111_011011_01010; 
		4965: oled_colour = 16'b01011_010100_01000; 
		4966: oled_colour = 16'b01111_011100_01011; 
		4967: oled_colour = 16'b10000_011110_01011; 
		4968: oled_colour = 16'b01001_010010_01000; 
		4969: oled_colour = 16'b01101_011000_01010; 
		4970: oled_colour = 16'b10001_100000_01011; 
		4971: oled_colour = 16'b01100_010101_01000; 
		4972: oled_colour = 16'b01101_011000_01001; 
		4973: oled_colour = 16'b10001_011111_01100; 
		4974: oled_colour = 16'b01100_010110_01001; 
		4975: oled_colour = 16'b01100_010110_01001; 
		4976: oled_colour = 16'b10000_011101_01011; 
		4977: oled_colour = 16'b01110_011001_01001; 
		4978: oled_colour = 16'b01100_010111_01001; 
		4979: oled_colour = 16'b10000_011110_01011; 
		4980: oled_colour = 16'b01110_011000_01001; 
		4981: oled_colour = 16'b01011_010101_01000; 
		4982: oled_colour = 16'b10001_100000_01100; 
		4983: oled_colour = 16'b01100_010110_01001; 
		4984: oled_colour = 16'b00111_001110_00111; 
		4985: oled_colour = 16'b01101_011000_01010; 
		4986: oled_colour = 16'b10001_100001_01100; 
		4987: oled_colour = 16'b10101_100111_01110; 
		4988: oled_colour = 16'b11010_110000_10000; 
		4989: oled_colour = 16'b11011_110010_10000; 
		4990: oled_colour = 16'b10100_100110_01101; 
		4991: oled_colour = 16'b01010_010010_01000; 
		4992: oled_colour = 16'b01111_010011_00010; 
		4993: oled_colour = 16'b01111_010101_00011; 
		4994: oled_colour = 16'b10001_010111_00011; 
		4995: oled_colour = 16'b10001_010111_00011; 
		4996: oled_colour = 16'b10001_010110_00011; 
		4997: oled_colour = 16'b10000_010101_00011; 
		4998: oled_colour = 16'b10000_010101_00011; 
		4999: oled_colour = 16'b10000_010101_00011; 
		5000: oled_colour = 16'b10001_010111_00100; 
		5001: oled_colour = 16'b10001_010111_00100; 
		5002: oled_colour = 16'b10001_010111_00100; 
		5003: oled_colour = 16'b10000_010110_00011; 
		5004: oled_colour = 16'b10000_010110_00011; 
		5005: oled_colour = 16'b10000_010110_00011; 
		5006: oled_colour = 16'b10000_010101_00011; 
		5007: oled_colour = 16'b10001_010111_00011; 
		5008: oled_colour = 16'b10001_011000_00100; 
		5009: oled_colour = 16'b10001_010111_00011; 
		5010: oled_colour = 16'b10000_010110_00011; 
		5011: oled_colour = 16'b10010_011010_00100; 
		5012: oled_colour = 16'b10000_010101_00011; 
		5013: oled_colour = 16'b10001_010111_00011; 
		5014: oled_colour = 16'b10000_010110_00011; 
		5015: oled_colour = 16'b10000_010110_00011; 
		5016: oled_colour = 16'b01111_010011_00010; 
		5017: oled_colour = 16'b01110_010011_00010; 
		5018: oled_colour = 16'b01111_010100_00010; 
		5019: oled_colour = 16'b10000_010110_00011; 
		5020: oled_colour = 16'b10001_010111_00011; 
		5021: oled_colour = 16'b01111_010100_00010; 
		5022: oled_colour = 16'b01111_010101_00011; 
		5023: oled_colour = 16'b10001_010111_00100; 
		5024: oled_colour = 16'b10010_011000_00100; 
		5025: oled_colour = 16'b10010_011001_00100; 
		5026: oled_colour = 16'b10000_010110_00011; 
		5027: oled_colour = 16'b10001_010110_00011; 
		5028: oled_colour = 16'b10000_010110_00011; 
		5029: oled_colour = 16'b10000_010101_00011; 
		5030: oled_colour = 16'b01111_010100_00010; 
		5031: oled_colour = 16'b10000_010110_00011; 
		5032: oled_colour = 16'b10010_011000_00100; 
		5033: oled_colour = 16'b10001_010111_00100; 
		5034: oled_colour = 16'b10001_010110_00011; 
		5035: oled_colour = 16'b10001_010111_00100; 
		5036: oled_colour = 16'b10001_010110_00011; 
		5037: oled_colour = 16'b10001_010111_00011; 
		5038: oled_colour = 16'b10010_011001_00100; 
		5039: oled_colour = 16'b10000_010101_00011; 
		5040: oled_colour = 16'b10010_011001_00101; 
		5041: oled_colour = 16'b10001_011000_00100; 
		5042: oled_colour = 16'b10000_010101_00011; 
		5043: oled_colour = 16'b01111_010101_00011; 
		5044: oled_colour = 16'b01111_010100_00011; 
		5045: oled_colour = 16'b10000_010110_00011; 
		5046: oled_colour = 16'b10000_010110_00011; 
		5047: oled_colour = 16'b10000_010101_00010; 
		5048: oled_colour = 16'b01111_010100_00010; 
		5049: oled_colour = 16'b10010_011000_00100; 
		5050: oled_colour = 16'b10011_011010_00100; 
		5051: oled_colour = 16'b10010_011001_00100; 
		5052: oled_colour = 16'b10011_011011_00101; 
		5053: oled_colour = 16'b10011_011011_00100; 
		5054: oled_colour = 16'b10011_011010_00100; 
		5055: oled_colour = 16'b10011_011010_00100; 
		5056: oled_colour = 16'b10001_010111_00100; 
		5057: oled_colour = 16'b10000_010110_00011; 
		5058: oled_colour = 16'b10010_011001_00100; 
		5059: oled_colour = 16'b10010_011000_00100; 
		5060: oled_colour = 16'b10010_011001_00100; 
		5061: oled_colour = 16'b10010_011001_00100; 
		5062: oled_colour = 16'b10011_011100_00101; 
		5063: oled_colour = 16'b10011_011011_00101; 
		5064: oled_colour = 16'b10010_011001_00100; 
		5065: oled_colour = 16'b10001_011000_00100; 
		5066: oled_colour = 16'b10001_011000_00011; 
		5067: oled_colour = 16'b10010_011010_00100; 
		5068: oled_colour = 16'b10011_011011_00100; 
		5069: oled_colour = 16'b10010_011001_00100; 
		5070: oled_colour = 16'b10010_011001_00100; 
		5071: oled_colour = 16'b10001_010111_00011; 
		5072: oled_colour = 16'b10001_010111_00100; 
		5073: oled_colour = 16'b10010_011010_00100; 
		5074: oled_colour = 16'b10010_011011_00100; 
		5075: oled_colour = 16'b10001_011000_00011; 
		5076: oled_colour = 16'b10011_011100_00101; 
		5077: oled_colour = 16'b10010_011011_00100; 
		5078: oled_colour = 16'b10011_011010_00100; 
		5079: oled_colour = 16'b10010_011000_00100; 
		5080: oled_colour = 16'b10001_011001_00100; 
		5081: oled_colour = 16'b10010_011010_00100; 
		5082: oled_colour = 16'b10010_011010_00100; 
		5083: oled_colour = 16'b10010_011001_00100; 
		5084: oled_colour = 16'b10010_011001_00100; 
		5085: oled_colour = 16'b10010_011001_00100; 
		5086: oled_colour = 16'b10010_011001_00100; 
		5087: oled_colour = 16'b10010_011001_00100; 
		5088: oled_colour = 16'b10011_011011_00101; 
		5089: oled_colour = 16'b10101_011110_00110; 
		5090: oled_colour = 16'b10011_011011_00101; 
		5091: oled_colour = 16'b10011_011011_00101; 
		5092: oled_colour = 16'b10011_011011_00101; 
		5093: oled_colour = 16'b10100_011101_00101; 
		5094: oled_colour = 16'b10100_011101_00101; 
		5095: oled_colour = 16'b10001_011000_00011; 
		5096: oled_colour = 16'b10011_011010_00101; 
		5097: oled_colour = 16'b10011_011011_00101; 
		5098: oled_colour = 16'b10011_011010_00101; 
		5099: oled_colour = 16'b10011_011010_00101; 
		5100: oled_colour = 16'b10011_011011_00101; 
		5101: oled_colour = 16'b10001_011000_00100; 
		5102: oled_colour = 16'b10100_011110_00110; 
		5103: oled_colour = 16'b10111_100011_01000; 
		5104: oled_colour = 16'b10011_011010_00100; 
		5105: oled_colour = 16'b10010_011001_00100; 
		5106: oled_colour = 16'b10010_011001_00100; 
		5107: oled_colour = 16'b10010_011001_00100; 
		5108: oled_colour = 16'b10010_011000_00100; 
		5109: oled_colour = 16'b10010_011010_00101; 
		5110: oled_colour = 16'b10010_011010_00100; 
		5111: oled_colour = 16'b10001_010111_00011; 
		5112: oled_colour = 16'b10011_011010_00101; 
		5113: oled_colour = 16'b10101_011111_00110; 
		5114: oled_colour = 16'b10011_011011_00100; 
		5115: oled_colour = 16'b10100_011101_00101; 
		5116: oled_colour = 16'b10010_011010_00100; 
		5117: oled_colour = 16'b10010_011001_00100; 
		5118: oled_colour = 16'b10011_011011_00101; 
		5119: oled_colour = 16'b10101_011110_00110; 
		5120: oled_colour = 16'b10011_011100_00101; 
		5121: oled_colour = 16'b10011_011100_00101; 
		5122: oled_colour = 16'b10011_011100_00101; 
		5123: oled_colour = 16'b10101_011111_00110; 
		5124: oled_colour = 16'b10101_011110_00110; 
		5125: oled_colour = 16'b10011_011011_00101; 
		5126: oled_colour = 16'b10001_011000_00100; 
		5127: oled_colour = 16'b10010_011010_00101; 
		5128: oled_colour = 16'b10100_011100_00110; 
		5129: oled_colour = 16'b10011_011011_00101; 
		5130: oled_colour = 16'b10011_011010_00101; 
		5131: oled_colour = 16'b10011_011010_00101; 
		5132: oled_colour = 16'b10010_011000_00100; 
		5133: oled_colour = 16'b10011_011001_00100; 
		5134: oled_colour = 16'b10011_011011_00101; 
		5135: oled_colour = 16'b10010_011001_00101; 
		5136: oled_colour = 16'b10101_011110_00110; 
		5137: oled_colour = 16'b10110_100000_00111; 
		5138: oled_colour = 16'b10101_011111_00110; 
		5139: oled_colour = 16'b10100_011101_00101; 
		5140: oled_colour = 16'b10001_010110_00011; 
		5141: oled_colour = 16'b10010_011001_00100; 
		5142: oled_colour = 16'b10010_011001_00100; 
		5143: oled_colour = 16'b10001_010111_00011; 
		5144: oled_colour = 16'b10010_011001_00100; 
		5145: oled_colour = 16'b10011_011010_00101; 
		5146: oled_colour = 16'b10011_011001_00101; 
		5147: oled_colour = 16'b10001_010111_00100; 
		5148: oled_colour = 16'b10010_011000_00100; 
		5149: oled_colour = 16'b10010_011001_00101; 
		5150: oled_colour = 16'b10011_011001_00101; 
		5151: oled_colour = 16'b10100_011100_00110; 
		5152: oled_colour = 16'b10011_011011_00101; 
		5153: oled_colour = 16'b10001_010111_00100; 
		5154: oled_colour = 16'b10010_011001_00101; 
		5155: oled_colour = 16'b10100_011100_00101; 
		5156: oled_colour = 16'b10101_011111_00111; 
		5157: oled_colour = 16'b10100_011101_00101; 
		5158: oled_colour = 16'b10011_011010_00101; 
		5159: oled_colour = 16'b10011_011011_00101; 
		5160: oled_colour = 16'b10100_011101_00110; 
		5161: oled_colour = 16'b10011_011100_00101; 
		5162: oled_colour = 16'b10001_011001_00100; 
		5163: oled_colour = 16'b10010_011001_00100; 
		5164: oled_colour = 16'b10011_011011_00101; 
		5165: oled_colour = 16'b10010_011010_00100; 
		5166: oled_colour = 16'b10011_011011_00101; 
		5167: oled_colour = 16'b10100_011100_00101; 
		5168: oled_colour = 16'b10001_010111_00011; 
		5169: oled_colour = 16'b10010_011000_00100; 
		5170: oled_colour = 16'b10010_011010_00101; 
		5171: oled_colour = 16'b10010_011001_00100; 
		5172: oled_colour = 16'b10001_011000_00100; 
		5173: oled_colour = 16'b10010_011000_00100; 
		5174: oled_colour = 16'b10010_011000_00100; 
		5175: oled_colour = 16'b10010_011000_00100; 
		5176: oled_colour = 16'b10101_100000_00111; 
		5177: oled_colour = 16'b10110_100001_00111; 
		5178: oled_colour = 16'b10001_011000_00100; 
		5179: oled_colour = 16'b10010_011010_00101; 
		5180: oled_colour = 16'b10011_011011_00101; 
		5181: oled_colour = 16'b10010_011001_00100; 
		5182: oled_colour = 16'b10011_011011_00101; 
		5183: oled_colour = 16'b10011_011001_00101; 
		5184: oled_colour = 16'b10100_011101_00110; 
		5185: oled_colour = 16'b10011_011010_00101; 
		5186: oled_colour = 16'b10011_011011_00101; 
		5187: oled_colour = 16'b10100_011111_00110; 
		5188: oled_colour = 16'b10101_011111_00110; 
		5189: oled_colour = 16'b10100_011101_00101; 
		5190: oled_colour = 16'b10010_011010_00100; 
		5191: oled_colour = 16'b10010_011001_00100; 
		5192: oled_colour = 16'b10010_011001_00100; 
		5193: oled_colour = 16'b10100_011101_00110; 
		5194: oled_colour = 16'b10010_011010_00101; 
		5195: oled_colour = 16'b10011_011011_00101; 
		5196: oled_colour = 16'b10101_100000_00110; 
		5197: oled_colour = 16'b10010_011001_00100; 
		5198: oled_colour = 16'b10110_100001_00111; 
		5199: oled_colour = 16'b10110_100000_00110; 
		5200: oled_colour = 16'b10010_011000_00100; 
		5201: oled_colour = 16'b10011_011001_00101; 
		5202: oled_colour = 16'b10011_011011_00101; 
		5203: oled_colour = 16'b10010_011000_00100; 
		5204: oled_colour = 16'b10011_011100_00101; 
		5205: oled_colour = 16'b10101_100000_00111; 
		5206: oled_colour = 16'b10011_011011_00101; 
		5207: oled_colour = 16'b10011_011010_00101; 
		5208: oled_colour = 16'b10101_011111_00111; 
		5209: oled_colour = 16'b10110_100010_00111; 
		5210: oled_colour = 16'b10111_100011_00111; 
		5211: oled_colour = 16'b10101_100001_00110; 
		5212: oled_colour = 16'b10001_010111_00100; 
		5213: oled_colour = 16'b10011_011101_00101; 
		5214: oled_colour = 16'b10011_011011_00101; 
		5215: oled_colour = 16'b10011_011010_00101; 
		5216: oled_colour = 16'b10110_100000_00111; 
		5217: oled_colour = 16'b10100_011110_00110; 
		5218: oled_colour = 16'b10101_011110_00110; 
		5219: oled_colour = 16'b10110_100001_00111; 
		5220: oled_colour = 16'b10100_011101_00110; 
		5221: oled_colour = 16'b10010_011001_00100; 
		5222: oled_colour = 16'b10011_011010_00101; 
		5223: oled_colour = 16'b10101_011111_00110; 
		5224: oled_colour = 16'b10101_011111_00111; 
		5225: oled_colour = 16'b10010_011010_00100; 
		5226: oled_colour = 16'b10010_011001_00101; 
		5227: oled_colour = 16'b10110_100000_00111; 
		5228: oled_colour = 16'b11000_100101_01000; 
		5229: oled_colour = 16'b11000_100110_01000; 
		5230: oled_colour = 16'b11000_100100_00111; 
		5231: oled_colour = 16'b10010_011001_00100; 
		5232: oled_colour = 16'b10100_011110_00110; 
		5233: oled_colour = 16'b10100_011101_00101; 
		5234: oled_colour = 16'b10100_011110_00101; 
		5235: oled_colour = 16'b11000_100100_01000; 
		5236: oled_colour = 16'b11000_100100_01000; 
		5237: oled_colour = 16'b10100_011101_00101; 
		5238: oled_colour = 16'b10010_011000_00100; 
		5239: oled_colour = 16'b10010_011001_00100; 
		5240: oled_colour = 16'b10011_011010_00101; 
		5241: oled_colour = 16'b10101_011111_00110; 
		5242: oled_colour = 16'b11001_100111_01001; 
		5243: oled_colour = 16'b11000_100101_01000; 
		5244: oled_colour = 16'b10111_100100_01000; 
		5245: oled_colour = 16'b10101_011110_00110; 
		5246: oled_colour = 16'b10010_011000_00100; 
		5247: oled_colour = 16'b10100_011100_00110; 
		5248: oled_colour = 16'b10101_011110_00111; 
		5249: oled_colour = 16'b10101_011111_00110; 
		5250: oled_colour = 16'b10010_011001_00100; 
		5251: oled_colour = 16'b10011_011010_00101; 
		5252: oled_colour = 16'b10101_011110_00110; 
		5253: oled_colour = 16'b10110_100001_00111; 
		5254: oled_colour = 16'b10100_011101_00101; 
		5255: oled_colour = 16'b10101_100000_00111; 
		5256: oled_colour = 16'b10101_011110_00110; 
		5257: oled_colour = 16'b10011_011011_00101; 
		5258: oled_colour = 16'b10011_011101_00101; 
		5259: oled_colour = 16'b10011_011011_00101; 
		5260: oled_colour = 16'b10010_011000_00100; 
		5261: oled_colour = 16'b10111_100100_01000; 
		5262: oled_colour = 16'b10111_100011_00111; 
		5263: oled_colour = 16'b10111_100010_00111; 
		5264: oled_colour = 16'b10100_011101_00110; 
		5265: oled_colour = 16'b10011_011010_00101; 
		5266: oled_colour = 16'b10100_011100_00101; 
		5267: oled_colour = 16'b10101_011111_00110; 
		5268: oled_colour = 16'b10010_011010_00100; 
		5269: oled_colour = 16'b10010_011001_00100; 
		5270: oled_colour = 16'b10011_011011_00101; 
		5271: oled_colour = 16'b10011_011001_00101; 
		5272: oled_colour = 16'b10010_011001_00100; 
		5273: oled_colour = 16'b10111_100011_01000; 
		5274: oled_colour = 16'b10100_011101_00110; 
		5275: oled_colour = 16'b10011_011100_00101; 
		5276: oled_colour = 16'b10101_011111_00110; 
		5277: oled_colour = 16'b10011_011010_00101; 
		5278: oled_colour = 16'b10011_011010_00101; 
		5279: oled_colour = 16'b10100_011100_00110; 
		5280: oled_colour = 16'b10100_011101_00101; 
		5281: oled_colour = 16'b10100_011101_00110; 
		5282: oled_colour = 16'b10100_011110_00110; 
		5283: oled_colour = 16'b10101_011111_00110; 
		5284: oled_colour = 16'b10100_011110_00110; 
		5285: oled_colour = 16'b10101_011111_00110; 
		5286: oled_colour = 16'b10110_100000_00111; 
		5287: oled_colour = 16'b10101_011111_00110; 
		5288: oled_colour = 16'b10110_100001_00111; 
		5289: oled_colour = 16'b10100_011110_00110; 
		5290: oled_colour = 16'b10100_011110_00110; 
		5291: oled_colour = 16'b11000_100110_01000; 
		5292: oled_colour = 16'b10101_100000_00110; 
		5293: oled_colour = 16'b10100_011101_00101; 
		5294: oled_colour = 16'b10101_011111_00110; 
		5295: oled_colour = 16'b10111_100011_00111; 
		5296: oled_colour = 16'b10101_011111_00110; 
		5297: oled_colour = 16'b10101_011111_00110; 
		5298: oled_colour = 16'b10100_011101_00110; 
		5299: oled_colour = 16'b10110_100001_00110; 
		5300: oled_colour = 16'b11000_100101_01000; 
		5301: oled_colour = 16'b10101_011111_00110; 
		5302: oled_colour = 16'b10100_011100_00101; 
		5303: oled_colour = 16'b10101_011111_00110; 
		5304: oled_colour = 16'b10101_100000_00110; 
		5305: oled_colour = 16'b10111_100100_00111; 
		5306: oled_colour = 16'b11001_100111_01000; 
		5307: oled_colour = 16'b10110_100010_00111; 
		5308: oled_colour = 16'b10101_011111_00110; 
		5309: oled_colour = 16'b10101_011110_00110; 
		5310: oled_colour = 16'b10101_100000_00110; 
		5311: oled_colour = 16'b10111_100011_01000; 
		5312: oled_colour = 16'b11000_100110_01000; 
		5313: oled_colour = 16'b10111_100100_00111; 
		5314: oled_colour = 16'b10111_100100_01000; 
		5315: oled_colour = 16'b10110_100010_00111; 
		5316: oled_colour = 16'b10011_011011_00101; 
		5317: oled_colour = 16'b10011_011100_00101; 
		5318: oled_colour = 16'b10101_100000_00110; 
		5319: oled_colour = 16'b10110_100010_00111; 
		5320: oled_colour = 16'b10110_100000_00110; 
		5321: oled_colour = 16'b10100_011101_00110; 
		5322: oled_colour = 16'b10101_011111_00110; 
		5323: oled_colour = 16'b11001_100111_01001; 
		5324: oled_colour = 16'b11001_100111_01000; 
		5325: oled_colour = 16'b11001_100111_01000; 
		5326: oled_colour = 16'b11001_100111_01000; 
		5327: oled_colour = 16'b10100_011110_00101; 
		5328: oled_colour = 16'b10101_011111_00110; 
		5329: oled_colour = 16'b10101_011111_00110; 
		5330: oled_colour = 16'b11010_101001_01001; 
		5331: oled_colour = 16'b11000_100101_01000; 
		5332: oled_colour = 16'b11000_100110_01000; 
		5333: oled_colour = 16'b11001_101000_01000; 
		5334: oled_colour = 16'b10011_011010_00101; 
		5335: oled_colour = 16'b10011_011011_00101; 
		5336: oled_colour = 16'b10011_011011_00101; 
		5337: oled_colour = 16'b10110_100001_00111; 
		5338: oled_colour = 16'b11010_101010_01001; 
		5339: oled_colour = 16'b11001_100111_01000; 
		5340: oled_colour = 16'b11001_101000_01001; 
		5341: oled_colour = 16'b11001_100111_01000; 
		5342: oled_colour = 16'b10101_011111_00110; 
		5343: oled_colour = 16'b10100_011101_00110; 
		5344: oled_colour = 16'b10110_100000_00111; 
		5345: oled_colour = 16'b10110_100010_00111; 
		5346: oled_colour = 16'b10101_100000_00110; 
		5347: oled_colour = 16'b10011_011011_00101; 
		5348: oled_colour = 16'b10100_011100_00101; 
		5349: oled_colour = 16'b10110_100010_00111; 
		5350: oled_colour = 16'b10111_100011_00111; 
		5351: oled_colour = 16'b11000_100100_01000; 
		5352: oled_colour = 16'b11001_100110_01000; 
		5353: oled_colour = 16'b10111_100011_00111; 
		5354: oled_colour = 16'b10101_011111_00110; 
		5355: oled_colour = 16'b10100_011110_00110; 
		5356: oled_colour = 16'b10101_100000_00110; 
		5357: oled_colour = 16'b10111_100011_00111; 
		5358: oled_colour = 16'b11000_100110_01000; 
		5359: oled_colour = 16'b10111_100100_00111; 
		5360: oled_colour = 16'b10110_100001_00110; 
		5361: oled_colour = 16'b10101_011110_00110; 
		5362: oled_colour = 16'b10100_011100_00101; 
		5363: oled_colour = 16'b10101_100000_00111; 
		5364: oled_colour = 16'b10111_100100_01000; 
		5365: oled_colour = 16'b10110_100001_00111; 
		5366: oled_colour = 16'b10100_011110_00110; 
		5367: oled_colour = 16'b10101_011110_00110; 
		5368: oled_colour = 16'b10101_011111_00110; 
		5369: oled_colour = 16'b10111_100010_00111; 
		5370: oled_colour = 16'b10101_011111_00110; 
		5371: oled_colour = 16'b10100_011101_00101; 
		5372: oled_colour = 16'b10110_100000_00111; 
		5373: oled_colour = 16'b11000_100101_01000; 
		5374: oled_colour = 16'b10101_011110_00101; 
		5375: oled_colour = 16'b10100_011101_00110; 
		5376: oled_colour = 16'b10101_011111_00110; 
		5377: oled_colour = 16'b10011_011011_00100; 
		5378: oled_colour = 16'b10010_011010_00100; 
		5379: oled_colour = 16'b10110_100000_00111; 
		5380: oled_colour = 16'b10110_100001_00111; 
		5381: oled_colour = 16'b10100_011101_00110; 
		5382: oled_colour = 16'b10110_100010_00111; 
		5383: oled_colour = 16'b10110_100000_00111; 
		5384: oled_colour = 16'b10011_011011_00101; 
		5385: oled_colour = 16'b10001_011000_00100; 
		5386: oled_colour = 16'b11000_100110_01000; 
		5387: oled_colour = 16'b11010_101010_01001; 
		5388: oled_colour = 16'b10100_011101_00101; 
		5389: oled_colour = 16'b11000_100100_01000; 
		5390: oled_colour = 16'b10111_100100_00111; 
		5391: oled_colour = 16'b10111_100100_01000; 
		5392: oled_colour = 16'b10101_011111_00110; 
		5393: oled_colour = 16'b10100_011110_00110; 
		5394: oled_colour = 16'b11001_101000_01000; 
		5395: oled_colour = 16'b11010_101011_01001; 
		5396: oled_colour = 16'b10111_100010_00111; 
		5397: oled_colour = 16'b10110_100010_00111; 
		5398: oled_colour = 16'b10101_100000_00110; 
		5399: oled_colour = 16'b10101_011110_00110; 
		5400: oled_colour = 16'b11010_101001_01001; 
		5401: oled_colour = 16'b11001_100111_01000; 
		5402: oled_colour = 16'b10110_100010_00111; 
		5403: oled_colour = 16'b10110_100011_00111; 
		5404: oled_colour = 16'b11001_100111_01000; 
		5405: oled_colour = 16'b10110_100001_00110; 
		5406: oled_colour = 16'b10101_100000_00110; 
		5407: oled_colour = 16'b11001_101000_01000; 
		5408: oled_colour = 16'b11010_101011_01001; 
		5409: oled_colour = 16'b10111_100100_01000; 
		5410: oled_colour = 16'b10110_100010_00111; 
		5411: oled_colour = 16'b10110_100010_00111; 
		5412: oled_colour = 16'b10111_100011_01000; 
		5413: oled_colour = 16'b10011_011011_00101; 
		5414: oled_colour = 16'b11000_100110_01000; 
		5415: oled_colour = 16'b11000_100110_01000; 
		5416: oled_colour = 16'b11010_101001_01001; 
		5417: oled_colour = 16'b10111_100100_00111; 
		5418: oled_colour = 16'b11000_100110_01000; 
		5419: oled_colour = 16'b11001_100111_01000; 
		5420: oled_colour = 16'b11001_100111_01000; 
		5421: oled_colour = 16'b11001_101000_01000; 
		5422: oled_colour = 16'b11000_100101_01000; 
		5423: oled_colour = 16'b10101_011111_00110; 
		5424: oled_colour = 16'b10111_100011_00111; 
		5425: oled_colour = 16'b10110_100010_00111; 
		5426: oled_colour = 16'b11001_101000_01000; 
		5427: oled_colour = 16'b11000_100110_01000; 
		5428: oled_colour = 16'b11000_100110_01000; 
		5429: oled_colour = 16'b11010_101011_01010; 
		5430: oled_colour = 16'b10100_011101_00101; 
		5431: oled_colour = 16'b10101_011110_00110; 
		5432: oled_colour = 16'b10110_100000_00111; 
		5433: oled_colour = 16'b10101_011111_00110; 
		5434: oled_colour = 16'b10110_100010_00111; 
		5435: oled_colour = 16'b11001_101000_01001; 
		5436: oled_colour = 16'b11001_100111_01000; 
		5437: oled_colour = 16'b11001_100111_01000; 
		5438: oled_colour = 16'b11001_100111_01000; 
		5439: oled_colour = 16'b10111_100010_00111; 
		5440: oled_colour = 16'b11010_101001_01001; 
		5441: oled_colour = 16'b11000_100110_01000; 
		5442: oled_colour = 16'b11001_101000_01001; 
		5443: oled_colour = 16'b10100_011101_00101; 
		5444: oled_colour = 16'b10110_100000_00111; 
		5445: oled_colour = 16'b10110_100010_00111; 
		5446: oled_colour = 16'b10111_100011_00111; 
		5447: oled_colour = 16'b10111_100011_00111; 
		5448: oled_colour = 16'b11010_101001_01001; 
		5449: oled_colour = 16'b11010_101010_01001; 
		5450: oled_colour = 16'b10110_100010_00111; 
		5451: oled_colour = 16'b10101_100000_00110; 
		5452: oled_colour = 16'b11000_100101_01000; 
		5453: oled_colour = 16'b10111_100100_00111; 
		5454: oled_colour = 16'b10101_100001_00110; 
		5455: oled_colour = 16'b11000_100110_01000; 
		5456: oled_colour = 16'b11001_101000_01001; 
		5457: oled_colour = 16'b10110_100010_00111; 
		5458: oled_colour = 16'b10101_011110_00110; 
		5459: oled_colour = 16'b10111_100010_00111; 
		5460: oled_colour = 16'b10110_100010_00111; 
		5461: oled_colour = 16'b11001_101000_01001; 
		5462: oled_colour = 16'b11010_101001_01000; 
		5463: oled_colour = 16'b10110_100010_00110; 
		5464: oled_colour = 16'b10100_011101_00110; 
		5465: oled_colour = 16'b10111_100100_01000; 
		5466: oled_colour = 16'b10111_100011_00111; 
		5467: oled_colour = 16'b11000_100110_01000; 
		5468: oled_colour = 16'b10100_011101_00101; 
		5469: oled_colour = 16'b11001_100111_01000; 
		5470: oled_colour = 16'b11001_101001_01001; 
		5471: oled_colour = 16'b10011_011100_00101; 
		5472: oled_colour = 16'b10110_100010_00111; 
		5473: oled_colour = 16'b10100_011110_00110; 
		5474: oled_colour = 16'b10110_100010_00111; 
		5475: oled_colour = 16'b11000_100110_01000; 
		5476: oled_colour = 16'b10101_011110_00110; 
		5477: oled_colour = 16'b10110_100000_00111; 
		5478: oled_colour = 16'b10101_011111_00110; 
		5479: oled_colour = 16'b10001_010111_00100; 
		5480: oled_colour = 16'b10010_011001_00100; 
		5481: oled_colour = 16'b10111_100100_00111; 
		5482: oled_colour = 16'b11010_101010_01001; 
		5483: oled_colour = 16'b11010_101010_01001; 
		5484: oled_colour = 16'b10100_011101_00101; 
		5485: oled_colour = 16'b10100_011101_00101; 
		5486: oled_colour = 16'b11011_101101_01010; 
		5487: oled_colour = 16'b11000_100101_01000; 
		5488: oled_colour = 16'b10011_011010_00100; 
		5489: oled_colour = 16'b10111_100011_00111; 
		5490: oled_colour = 16'b10111_100100_00111; 
		5491: oled_colour = 16'b10110_100000_00110; 
		5492: oled_colour = 16'b10110_100001_00111; 
		5493: oled_colour = 16'b11000_100110_01000; 
		5494: oled_colour = 16'b11000_100101_01000; 
		5495: oled_colour = 16'b10111_100011_00111; 
		5496: oled_colour = 16'b11001_100111_01000; 
		5497: oled_colour = 16'b11001_100111_01000; 
		5498: oled_colour = 16'b10101_011111_00110; 
		5499: oled_colour = 16'b10110_100001_00110; 
		5500: oled_colour = 16'b10110_100010_00111; 
		5501: oled_colour = 16'b10111_100100_00111; 
		5502: oled_colour = 16'b11001_101000_01001; 
		5503: oled_colour = 16'b11001_101000_01001; 
		5504: oled_colour = 16'b11001_100111_01000; 
		5505: oled_colour = 16'b10101_011111_00110; 
		5506: oled_colour = 16'b10111_100101_01000; 
		5507: oled_colour = 16'b11001_101000_01001; 
		5508: oled_colour = 16'b10110_100010_00111; 
		5509: oled_colour = 16'b10101_100001_00110; 
		5510: oled_colour = 16'b11001_100111_01000; 
		5511: oled_colour = 16'b11001_101000_01000; 
		5512: oled_colour = 16'b11001_101000_01001; 
		5513: oled_colour = 16'b10101_100000_00110; 
		5514: oled_colour = 16'b11010_101001_01001; 
		5515: oled_colour = 16'b11001_101000_01000; 
		5516: oled_colour = 16'b11000_100101_00111; 
		5517: oled_colour = 16'b11000_100101_01000; 
		5518: oled_colour = 16'b10101_011111_00110; 
		5519: oled_colour = 16'b10101_011111_00110; 
		5520: oled_colour = 16'b10101_011110_00110; 
		5521: oled_colour = 16'b10100_011110_00110; 
		5522: oled_colour = 16'b10111_100100_00111; 
		5523: oled_colour = 16'b11010_101001_01000; 
		5524: oled_colour = 16'b11011_101011_01001; 
		5525: oled_colour = 16'b10110_100010_00111; 
		5526: oled_colour = 16'b10111_100011_00111; 
		5527: oled_colour = 16'b10110_100000_00111; 
		5528: oled_colour = 16'b10111_100010_00111; 
		5529: oled_colour = 16'b10111_100011_00111; 
		5530: oled_colour = 16'b10100_011101_00110; 
		5531: oled_colour = 16'b10110_100010_00111; 
		5532: oled_colour = 16'b11000_100101_00111; 
		5533: oled_colour = 16'b11000_100110_01000; 
		5534: oled_colour = 16'b11010_101001_01001; 
		5535: oled_colour = 16'b11000_100101_01000; 
		5536: oled_colour = 16'b10110_100010_00111; 
		5537: oled_colour = 16'b11010_101001_01001; 
		5538: oled_colour = 16'b11001_101000_01001; 
		5539: oled_colour = 16'b10111_100100_00111; 
		5540: oled_colour = 16'b10110_100000_00110; 
		5541: oled_colour = 16'b11000_100110_01000; 
		5542: oled_colour = 16'b11001_101000_01000; 
		5543: oled_colour = 16'b10110_100001_00111; 
		5544: oled_colour = 16'b10111_100010_00111; 
		5545: oled_colour = 16'b11001_101001_01001; 
		5546: oled_colour = 16'b11001_101000_01000; 
		5547: oled_colour = 16'b11000_100110_01000; 
		5548: oled_colour = 16'b10110_100011_00111; 
		5549: oled_colour = 16'b10110_100010_00111; 
		5550: oled_colour = 16'b10101_100001_00110; 
		5551: oled_colour = 16'b10110_100011_00111; 
		5552: oled_colour = 16'b11001_101000_01001; 
		5553: oled_colour = 16'b11000_100110_01000; 
		5554: oled_colour = 16'b10111_100010_00111; 
		5555: oled_colour = 16'b11001_100111_01000; 
		5556: oled_colour = 16'b10111_100011_00111; 
		5557: oled_colour = 16'b10110_100001_00111; 
		5558: oled_colour = 16'b10110_100010_00111; 
		5559: oled_colour = 16'b10111_100100_00111; 
		5560: oled_colour = 16'b10101_011110_00110; 
		5561: oled_colour = 16'b10100_011101_00101; 
		5562: oled_colour = 16'b11010_101010_01001; 
		5563: oled_colour = 16'b11001_101001_01000; 
		5564: oled_colour = 16'b10001_011000_00011; 
		5565: oled_colour = 16'b11000_100101_01000; 
		5566: oled_colour = 16'b11011_101011_01001; 
		5567: oled_colour = 16'b11010_101001_01001; 
		5568: oled_colour = 16'b11011_101100_01010; 
		5569: oled_colour = 16'b11001_100111_01000; 
		5570: oled_colour = 16'b11010_101010_01001; 
		5571: oled_colour = 16'b11010_101011_01001; 
		5572: oled_colour = 16'b10110_100010_00111; 
		5573: oled_colour = 16'b10101_100000_00110; 
		5574: oled_colour = 16'b10110_100010_00111; 
		5575: oled_colour = 16'b10111_100100_01000; 
		5576: oled_colour = 16'b11001_100111_01001; 
		5577: oled_colour = 16'b11011_101100_01010; 
		5578: oled_colour = 16'b11011_101100_01001; 
		5579: oled_colour = 16'b11000_100110_01000; 
		5580: oled_colour = 16'b10100_011101_00101; 
		5581: oled_colour = 16'b10110_100001_00110; 
		5582: oled_colour = 16'b11011_101101_01010; 
		5583: oled_colour = 16'b10110_100010_00110; 
		5584: oled_colour = 16'b11000_100101_01000; 
		5585: oled_colour = 16'b11010_101001_01001; 
		5586: oled_colour = 16'b10110_100001_00110; 
		5587: oled_colour = 16'b11010_101010_01001; 
		5588: oled_colour = 16'b11001_101000_01000; 
		5589: oled_colour = 16'b11000_100101_00111; 
		5590: oled_colour = 16'b11000_100110_01000; 
		5591: oled_colour = 16'b11001_100111_01000; 
		5592: oled_colour = 16'b11000_100110_01000; 
		5593: oled_colour = 16'b10111_100011_00111; 
		5594: oled_colour = 16'b11000_100110_01000; 
		5595: oled_colour = 16'b11001_101000_01001; 
		5596: oled_colour = 16'b11001_101000_01001; 
		5597: oled_colour = 16'b11001_101000_01001; 
		5598: oled_colour = 16'b11001_101000_01000; 
		5599: oled_colour = 16'b11010_101011_01001; 
		5600: oled_colour = 16'b11010_101001_01000; 
		5601: oled_colour = 16'b11001_100111_01000; 
		5602: oled_colour = 16'b11001_100111_01000; 
		5603: oled_colour = 16'b11011_101100_01010; 
		5604: oled_colour = 16'b10110_100011_00110; 
		5605: oled_colour = 16'b11001_101001_01001; 
		5606: oled_colour = 16'b11001_101000_01000; 
		5607: oled_colour = 16'b11001_101000_01000; 
		5608: oled_colour = 16'b10111_100011_00111; 
		5609: oled_colour = 16'b10111_100100_01000; 
		5610: oled_colour = 16'b11001_101000_01000; 
		5611: oled_colour = 16'b11001_100111_01000; 
		5612: oled_colour = 16'b10111_100100_00111; 
		5613: oled_colour = 16'b11000_100110_01000; 
		5614: oled_colour = 16'b10101_100000_00110; 
		5615: oled_colour = 16'b10110_100001_00110; 
		5616: oled_colour = 16'b11000_100101_00111; 
		5617: oled_colour = 16'b11000_100111_01000; 
		5618: oled_colour = 16'b11010_101011_01001; 
		5619: oled_colour = 16'b11011_101100_01010; 
		5620: oled_colour = 16'b10110_100001_00111; 
		5621: oled_colour = 16'b10011_011011_00101; 
		5622: oled_colour = 16'b10111_100011_01000; 
		5623: oled_colour = 16'b10110_100001_00111; 
		5624: oled_colour = 16'b10110_100010_00111; 
		5625: oled_colour = 16'b11010_101001_01001; 
		5626: oled_colour = 16'b10110_100001_00110; 
		5627: oled_colour = 16'b10110_100001_00111; 
		5628: oled_colour = 16'b11000_100101_00111; 
		5629: oled_colour = 16'b10111_100101_00111; 
		5630: oled_colour = 16'b11001_100111_01000; 
		5631: oled_colour = 16'b11001_100111_01000; 
		5632: oled_colour = 16'b10111_100100_01000; 
		5633: oled_colour = 16'b11000_100101_01000; 
		5634: oled_colour = 16'b11001_100111_01000; 
		5635: oled_colour = 16'b11010_101001_01001; 
		5636: oled_colour = 16'b11001_101000_01000; 
		5637: oled_colour = 16'b10111_100100_00111; 
		5638: oled_colour = 16'b11011_101100_01010; 
		5639: oled_colour = 16'b11000_100110_01000; 
		5640: oled_colour = 16'b11001_100111_01000; 
		5641: oled_colour = 16'b11010_101010_01001; 
		5642: oled_colour = 16'b11010_101010_01001; 
		5643: oled_colour = 16'b11010_101001_01001; 
		5644: oled_colour = 16'b11001_101000_01000; 
		5645: oled_colour = 16'b11001_101000_01001; 
		5646: oled_colour = 16'b11001_100111_01000; 
		5647: oled_colour = 16'b11000_100101_01000; 
		5648: oled_colour = 16'b10111_100100_00111; 
		5649: oled_colour = 16'b10111_100101_01000; 
		5650: oled_colour = 16'b11001_101000_01001; 
		5651: oled_colour = 16'b11000_100110_01000; 
		5652: oled_colour = 16'b11000_100101_00111; 
		5653: oled_colour = 16'b11001_101000_01000; 
		5654: oled_colour = 16'b11001_101001_01001; 
		5655: oled_colour = 16'b10111_100010_00110; 
		5656: oled_colour = 16'b11010_101001_01001; 
		5657: oled_colour = 16'b10111_100100_00111; 
		5658: oled_colour = 16'b11000_100101_00111; 
		5659: oled_colour = 16'b11011_101100_01010; 
		5660: oled_colour = 16'b10101_011111_00110; 
		5661: oled_colour = 16'b10101_011111_00110; 
		5662: oled_colour = 16'b11000_100110_01000; 
		5663: oled_colour = 16'b11011_101100_01010; 
		5664: oled_colour = 16'b11000_100110_01000; 
		5665: oled_colour = 16'b11000_100110_01000; 
		5666: oled_colour = 16'b11001_101000_01000; 
		5667: oled_colour = 16'b11000_100110_01000; 
		5668: oled_colour = 16'b11011_101100_01010; 
		5669: oled_colour = 16'b11011_101101_01010; 
		5670: oled_colour = 16'b11010_101011_01010; 
		5671: oled_colour = 16'b11010_101011_01001; 
		5672: oled_colour = 16'b11100_101110_01010; 
		5673: oled_colour = 16'b11100_101110_01010; 
		5674: oled_colour = 16'b10101_011111_00101; 
		5675: oled_colour = 16'b10011_011011_00100; 
		5676: oled_colour = 16'b11001_101000_01001; 
		5677: oled_colour = 16'b11000_100110_01000; 
		5678: oled_colour = 16'b11001_101000_01000; 
		5679: oled_colour = 16'b11011_101101_01010; 
		5680: oled_colour = 16'b11011_101011_01001; 
		5681: oled_colour = 16'b11001_100111_01000; 
		5682: oled_colour = 16'b11010_101001_01001; 
		5683: oled_colour = 16'b10111_100100_00111; 
		5684: oled_colour = 16'b10011_011100_00101; 
		5685: oled_colour = 16'b11010_101011_01001; 
		5686: oled_colour = 16'b11100_110000_01011; 
		5687: oled_colour = 16'b11000_100110_01000; 
		5688: oled_colour = 16'b10100_011111_00101; 
		5689: oled_colour = 16'b10111_100100_00111; 
		5690: oled_colour = 16'b11000_100101_01000; 
		5691: oled_colour = 16'b10111_100100_00111; 
		5692: oled_colour = 16'b11010_101001_01001; 
		5693: oled_colour = 16'b11010_101010_01001; 
		5694: oled_colour = 16'b11001_101000_01001; 
		5695: oled_colour = 16'b11000_100101_00111; 
		5696: oled_colour = 16'b11011_101011_01001; 
		5697: oled_colour = 16'b11001_101000_01000; 
		5698: oled_colour = 16'b11000_100110_01000; 
		5699: oled_colour = 16'b11010_101011_01010; 
		5700: oled_colour = 16'b11001_101000_01000; 
		5701: oled_colour = 16'b11011_101101_01010; 
		5702: oled_colour = 16'b11000_100101_01000; 
		5703: oled_colour = 16'b11000_100110_01000; 
		5704: oled_colour = 16'b11011_101100_01010; 
		5705: oled_colour = 16'b10111_100100_00111; 
		5706: oled_colour = 16'b10100_011101_00101; 
		5707: oled_colour = 16'b11010_101010_01001; 
		5708: oled_colour = 16'b10011_011100_00101; 
		5709: oled_colour = 16'b11001_100111_01000; 
		5710: oled_colour = 16'b10110_100010_00111; 
		5711: oled_colour = 16'b11001_101001_01001; 
		5712: oled_colour = 16'b11000_100110_01000; 
		5713: oled_colour = 16'b10101_011111_00110; 
		5714: oled_colour = 16'b11101_110001_01011; 
		5715: oled_colour = 16'b11001_100111_01000; 
		5716: oled_colour = 16'b10010_011000_00100; 
		5717: oled_colour = 16'b10000_010101_00010; 
		5718: oled_colour = 16'b10101_011111_00110; 
		5719: oled_colour = 16'b11000_100110_01000; 
		5720: oled_colour = 16'b11011_101011_01001; 
		5721: oled_colour = 16'b11011_101011_01010; 
		5722: oled_colour = 16'b11000_100111_01000; 
		5723: oled_colour = 16'b10101_100000_00110; 
		5724: oled_colour = 16'b11010_101010_01001; 
		5725: oled_colour = 16'b10010_011011_00100; 
		5726: oled_colour = 16'b11001_101001_01001; 
		5727: oled_colour = 16'b10101_100000_00110; 
		5728: oled_colour = 16'b10110_100010_00110; 
		5729: oled_colour = 16'b11010_101001_01001; 
		5730: oled_colour = 16'b11010_101001_01001; 
		5731: oled_colour = 16'b10111_100100_00111; 
		5732: oled_colour = 16'b11011_101100_01010; 
		5733: oled_colour = 16'b11001_101001_01001; 
		5734: oled_colour = 16'b11010_101010_01001; 
		5735: oled_colour = 16'b11001_101000_01000; 
		5736: oled_colour = 16'b11000_100110_01000; 
		5737: oled_colour = 16'b11010_101011_01001; 
		5738: oled_colour = 16'b11001_100111_01000; 
		5739: oled_colour = 16'b11000_100110_01000; 
		5740: oled_colour = 16'b11010_101010_01001; 
		5741: oled_colour = 16'b11010_101010_01001; 
		5742: oled_colour = 16'b11000_100101_01000; 
		5743: oled_colour = 16'b11000_100110_01000; 
		5744: oled_colour = 16'b10111_100100_00111; 
		5745: oled_colour = 16'b10101_100000_00110; 
		5746: oled_colour = 16'b10111_100011_00111; 
		5747: oled_colour = 16'b11100_101110_01010; 
		5748: oled_colour = 16'b11011_101101_01010; 
		5749: oled_colour = 16'b10101_100000_00110; 
		5750: oled_colour = 16'b10110_100001_00110; 
		5751: oled_colour = 16'b11001_101000_01001; 
		5752: oled_colour = 16'b11001_101000_01001; 
		5753: oled_colour = 16'b11010_101010_01001; 
		5754: oled_colour = 16'b11010_101011_01001; 
		5755: oled_colour = 16'b11010_101010_01001; 
		5756: oled_colour = 16'b11001_100111_01000; 
		5757: oled_colour = 16'b11000_100111_01000; 
		5758: oled_colour = 16'b10100_011110_00101; 
		5759: oled_colour = 16'b10011_011101_00101; 
		5760: oled_colour = 16'b11000_100101_00111; 
		5761: oled_colour = 16'b10101_100000_00110; 
		5762: oled_colour = 16'b10111_100011_00111; 
		5763: oled_colour = 16'b11000_100110_01000; 
		5764: oled_colour = 16'b11001_100111_01000; 
		5765: oled_colour = 16'b11001_100111_01000; 
		5766: oled_colour = 16'b11001_101000_01000; 
		5767: oled_colour = 16'b10111_100101_01000; 
		5768: oled_colour = 16'b10011_011100_00101; 
		5769: oled_colour = 16'b10000_010101_00010; 
		5770: oled_colour = 16'b10010_011010_00100; 
		5771: oled_colour = 16'b10110_100001_00110; 
		5772: oled_colour = 16'b11000_100101_00111; 
		5773: oled_colour = 16'b11001_101000_01000; 
		5774: oled_colour = 16'b11010_101001_01001; 
		5775: oled_colour = 16'b11000_100100_00111; 
		5776: oled_colour = 16'b10111_100100_00111; 
		5777: oled_colour = 16'b11010_101100_01010; 
		5778: oled_colour = 16'b10100_011111_00101; 
		5779: oled_colour = 16'b10001_010110_00011; 
		5780: oled_colour = 16'b11010_101011_01001; 
		5781: oled_colour = 16'b11100_101110_01010; 
		5782: oled_colour = 16'b10101_100000_00110; 
		5783: oled_colour = 16'b10011_011011_00100; 
		5784: oled_colour = 16'b11001_101001_01001; 
		5785: oled_colour = 16'b11010_101001_01001; 
		5786: oled_colour = 16'b11010_101010_01001; 
		5787: oled_colour = 16'b11100_110000_01011; 
		5788: oled_colour = 16'b11010_101010_01001; 
		5789: oled_colour = 16'b11001_101001_01001; 
		5790: oled_colour = 16'b10001_011000_00100; 
		5791: oled_colour = 16'b10111_100011_00111; 
		5792: oled_colour = 16'b10111_100011_00111; 
		5793: oled_colour = 16'b11000_100101_01000; 
		5794: oled_colour = 16'b11011_101100_01001; 
		5795: oled_colour = 16'b11001_101001_01000; 
		5796: oled_colour = 16'b11010_101011_01001; 
		5797: oled_colour = 16'b11010_101001_01001; 
		5798: oled_colour = 16'b11001_101001_01000; 
		5799: oled_colour = 16'b11101_110001_01010; 
		5800: oled_colour = 16'b10011_011011_00100; 
		5801: oled_colour = 16'b10010_011001_00101; 
		5802: oled_colour = 16'b11000_100110_01000; 
		5803: oled_colour = 16'b11000_100111_01000; 
		5804: oled_colour = 16'b10010_011001_00100; 
		5805: oled_colour = 16'b11010_101001_01001; 
		5806: oled_colour = 16'b10101_011111_00101; 
		5807: oled_colour = 16'b10010_011011_00101; 
		5808: oled_colour = 16'b10000_010100_00010; 
		5809: oled_colour = 16'b11010_101010_01001; 
		5810: oled_colour = 16'b11101_110000_01010; 
		5811: oled_colour = 16'b11001_100111_01000; 
		5812: oled_colour = 16'b10100_011100_00101; 
		5813: oled_colour = 16'b10001_010110_00011; 
		5814: oled_colour = 16'b10111_100011_00111; 
		5815: oled_colour = 16'b11010_101010_01001; 
		5816: oled_colour = 16'b10100_011101_00101; 
		5817: oled_colour = 16'b10111_100011_00111; 
		5818: oled_colour = 16'b11010_101011_01001; 
		5819: oled_colour = 16'b10100_011110_00101; 
		5820: oled_colour = 16'b11000_100101_01000; 
		5821: oled_colour = 16'b10110_100010_00110; 
		5822: oled_colour = 16'b10100_011101_00101; 
		5823: oled_colour = 16'b11010_101010_01001; 
		5824: oled_colour = 16'b10101_011110_00110; 
		5825: oled_colour = 16'b10010_011001_00100; 
		5826: oled_colour = 16'b11000_100110_01000; 
		5827: oled_colour = 16'b11100_101111_01010; 
		5828: oled_colour = 16'b11000_100110_01000; 
		5829: oled_colour = 16'b11011_101100_01010; 
		5830: oled_colour = 16'b11001_101001_01000; 
		5831: oled_colour = 16'b11010_101010_01001; 
		5832: oled_colour = 16'b11010_101010_01001; 
		5833: oled_colour = 16'b10110_100010_00110; 
		5834: oled_colour = 16'b11000_100110_01000; 
		5835: oled_colour = 16'b10011_011100_00100; 
		5836: oled_colour = 16'b10101_100001_00110; 
		5837: oled_colour = 16'b11010_101010_01001; 
		5838: oled_colour = 16'b11011_101101_01010; 
		5839: oled_colour = 16'b11100_101110_01010; 
		5840: oled_colour = 16'b11001_101001_01000; 
		5841: oled_colour = 16'b11010_101010_01001; 
		5842: oled_colour = 16'b10110_100010_00110; 
		5843: oled_colour = 16'b10011_011011_00100; 
		5844: oled_colour = 16'b11001_101000_01000; 
		5845: oled_colour = 16'b11100_101110_01010; 
		5846: oled_colour = 16'b10101_011111_00101; 
		5847: oled_colour = 16'b10010_011001_00100; 
		5848: oled_colour = 16'b11000_100110_01000; 
		5849: oled_colour = 16'b11010_101010_01001; 
		5850: oled_colour = 16'b10111_100100_00111; 
		5851: oled_colour = 16'b11001_100111_01000; 
		5852: oled_colour = 16'b11001_101000_01000; 
		5853: oled_colour = 16'b11001_100111_01000; 
		5854: oled_colour = 16'b10111_100011_00111; 
		5855: oled_colour = 16'b10011_011100_00101; 
		5856: oled_colour = 16'b11011_101101_01011; 
		5857: oled_colour = 16'b11010_101100_01011; 
		5858: oled_colour = 16'b11011_101111_01100; 
		5859: oled_colour = 16'b11100_110001_01101; 
		5860: oled_colour = 16'b11011_101110_01011; 
		5861: oled_colour = 16'b11011_101100_01010; 
		5862: oled_colour = 16'b10111_100011_00111; 
		5863: oled_colour = 16'b10010_011011_00101; 
		5864: oled_colour = 16'b10100_011110_00110; 
		5865: oled_colour = 16'b11001_101010_01011; 
		5866: oled_colour = 16'b11101_110011_01101; 
		5867: oled_colour = 16'b11000_101001_01010; 
		5868: oled_colour = 16'b11101_110001_01101; 
		5869: oled_colour = 16'b11101_110001_01100; 
		5870: oled_colour = 16'b11010_101011_01010; 
		5871: oled_colour = 16'b11001_101001_01010; 
		5872: oled_colour = 16'b11111_110110_01110; 
		5873: oled_colour = 16'b11010_101100_01010; 
		5874: oled_colour = 16'b10100_011110_00110; 
		5875: oled_colour = 16'b11001_101000_01010; 
		5876: oled_colour = 16'b11110_110101_01110; 
		5877: oled_colour = 16'b11101_110011_01101; 
		5878: oled_colour = 16'b11000_100111_01000; 
		5879: oled_colour = 16'b11011_101110_01100; 
		5880: oled_colour = 16'b11101_110011_01101; 
		5881: oled_colour = 16'b11011_101110_01010; 
		5882: oled_colour = 16'b11101_110011_01110; 
		5883: oled_colour = 16'b11110_110110_01110; 
		5884: oled_colour = 16'b11100_110000_01100; 
		5885: oled_colour = 16'b10111_100101_01000; 
		5886: oled_colour = 16'b10101_100000_00110; 
		5887: oled_colour = 16'b11101_110001_01101; 
		5888: oled_colour = 16'b10111_100100_00111; 
		5889: oled_colour = 16'b11100_101111_01100; 
		5890: oled_colour = 16'b11100_110001_01100; 
		5891: oled_colour = 16'b11011_101110_01011; 
		5892: oled_colour = 16'b11110_110100_01110; 
		5893: oled_colour = 16'b11011_101100_01010; 
		5894: oled_colour = 16'b11101_110010_01101; 
		5895: oled_colour = 16'b11110_110101_01110; 
		5896: oled_colour = 16'b11000_100111_01001; 
		5897: oled_colour = 16'b10111_100011_01000; 
		5898: oled_colour = 16'b11101_110001_01100; 
		5899: oled_colour = 16'b11001_101000_01001; 
		5900: oled_colour = 16'b11001_101001_01001; 
		5901: oled_colour = 16'b11101_110011_01101; 
		5902: oled_colour = 16'b10111_100110_01001; 
		5903: oled_colour = 16'b10101_100001_00110; 
		5904: oled_colour = 16'b11010_101101_01011; 
		5905: oled_colour = 16'b11111_111000_01111; 
		5906: oled_colour = 16'b11110_110101_01101; 
		5907: oled_colour = 16'b11101_110011_01101; 
		5908: oled_colour = 16'b11100_110000_01101; 
		5909: oled_colour = 16'b11001_101010_01010; 
		5910: oled_colour = 16'b11101_110001_01101; 
		5911: oled_colour = 16'b11101_110001_01101; 
		5912: oled_colour = 16'b10110_100100_00111; 
		5913: oled_colour = 16'b10111_100110_01000; 
		5914: oled_colour = 16'b11110_110100_01110; 
		5915: oled_colour = 16'b11010_101100_01011; 
		5916: oled_colour = 16'b11000_100111_01001; 
		5917: oled_colour = 16'b11110_110101_01110; 
		5918: oled_colour = 16'b10111_100101_01000; 
		5919: oled_colour = 16'b11011_101101_01011; 
		5920: oled_colour = 16'b11011_101110_01011; 
		5921: oled_colour = 16'b10101_100001_00111; 
		5922: oled_colour = 16'b11001_101011_01010; 
		5923: oled_colour = 16'b11111_111000_01111; 
		5924: oled_colour = 16'b11100_101111_01011; 
		5925: oled_colour = 16'b11100_101110_01011; 
		5926: oled_colour = 16'b11101_110011_01110; 
		5927: oled_colour = 16'b11011_101111_01100; 
		5928: oled_colour = 16'b11101_110010_01100; 
		5929: oled_colour = 16'b11010_101011_01010; 
		5930: oled_colour = 16'b11000_100111_01001; 
		5931: oled_colour = 16'b11100_101111_01100; 
		5932: oled_colour = 16'b10100_011110_00101; 
		5933: oled_colour = 16'b11001_101010_01010; 
		5934: oled_colour = 16'b11100_110000_01100; 
		5935: oled_colour = 16'b11111_110111_01111; 
		5936: oled_colour = 16'b11100_110001_01101; 
		5937: oled_colour = 16'b11100_101111_01011; 
		5938: oled_colour = 16'b11110_110011_01101; 
		5939: oled_colour = 16'b11001_101001_01010; 
		5940: oled_colour = 16'b11001_101001_01001; 
		5941: oled_colour = 16'b11111_110110_01110; 
		5942: oled_colour = 16'b11101_110010_01101; 
		5943: oled_colour = 16'b10110_100100_01000; 
		5944: oled_colour = 16'b10101_100000_00110; 
		5945: oled_colour = 16'b11101_110001_01100; 
		5946: oled_colour = 16'b11101_110010_01101; 
		5947: oled_colour = 16'b11001_101001_01010; 
		5948: oled_colour = 16'b11011_101101_01011; 
		5949: oled_colour = 16'b11101_110010_01101; 
		5950: oled_colour = 16'b11100_110000_01100; 
		5951: oled_colour = 16'b11010_101011_01010; 
		5952: oled_colour = 16'b11011_101100_01011; 
		5953: oled_colour = 16'b11011_101110_01011; 
		5954: oled_colour = 16'b11011_101110_01011; 
		5955: oled_colour = 16'b11011_101110_01011; 
		5956: oled_colour = 16'b11011_101101_01011; 
		5957: oled_colour = 16'b11100_101101_01010; 
		5958: oled_colour = 16'b10110_100001_00111; 
		5959: oled_colour = 16'b11000_100110_01000; 
		5960: oled_colour = 16'b11100_101111_01011; 
		5961: oled_colour = 16'b11100_101111_01011; 
		5962: oled_colour = 16'b11010_101100_01010; 
		5963: oled_colour = 16'b11001_101001_01010; 
		5964: oled_colour = 16'b11011_101110_01011; 
		5965: oled_colour = 16'b11011_101100_01011; 
		5966: oled_colour = 16'b11001_101001_01001; 
		5967: oled_colour = 16'b11011_101101_01011; 
		5968: oled_colour = 16'b11011_101110_01011; 
		5969: oled_colour = 16'b10110_100011_00111; 
		5970: oled_colour = 16'b11010_101001_01001; 
		5971: oled_colour = 16'b11100_101110_01011; 
		5972: oled_colour = 16'b11011_101100_01010; 
		5973: oled_colour = 16'b11011_101101_01011; 
		5974: oled_colour = 16'b11010_101011_01010; 
		5975: oled_colour = 16'b11100_101111_01100; 
		5976: oled_colour = 16'b11010_101011_01010; 
		5977: oled_colour = 16'b11010_101010_01001; 
		5978: oled_colour = 16'b11011_101101_01011; 
		5979: oled_colour = 16'b11011_101100_01011; 
		5980: oled_colour = 16'b11011_101110_01011; 
		5981: oled_colour = 16'b10111_100101_01000; 
		5982: oled_colour = 16'b11011_101100_01010; 
		5983: oled_colour = 16'b11011_101100_01011; 
		5984: oled_colour = 16'b11010_101010_01001; 
		5985: oled_colour = 16'b11011_101101_01011; 
		5986: oled_colour = 16'b11001_101010_01010; 
		5987: oled_colour = 16'b11010_101100_01011; 
		5988: oled_colour = 16'b11011_101110_01011; 
		5989: oled_colour = 16'b11010_101011_01010; 
		5990: oled_colour = 16'b11011_101100_01010; 
		5991: oled_colour = 16'b11011_101101_01011; 
		5992: oled_colour = 16'b11100_101111_01011; 
		5993: oled_colour = 16'b10111_100100_00111; 
		5994: oled_colour = 16'b11010_101010_01010; 
		5995: oled_colour = 16'b11000_100111_01000; 
		5996: oled_colour = 16'b11001_101000_01001; 
		5997: oled_colour = 16'b11100_101110_01011; 
		5998: oled_colour = 16'b11010_101010_01010; 
		5999: oled_colour = 16'b11000_100111_01000; 
		6000: oled_colour = 16'b11011_101110_01011; 
		6001: oled_colour = 16'b11011_101101_01011; 
		6002: oled_colour = 16'b11011_101100_01010; 
		6003: oled_colour = 16'b11011_101101_01011; 
		6004: oled_colour = 16'b11011_101101_01011; 
		6005: oled_colour = 16'b11100_101110_01011; 
		6006: oled_colour = 16'b11011_101101_01011; 
		6007: oled_colour = 16'b11011_101101_01011; 
		6008: oled_colour = 16'b11011_101011_01010; 
		6009: oled_colour = 16'b11100_101111_01011; 
		6010: oled_colour = 16'b11100_101111_01100; 
		6011: oled_colour = 16'b11010_101011_01010; 
		6012: oled_colour = 16'b11010_101011_01010; 
		6013: oled_colour = 16'b11100_101111_01011; 
		6014: oled_colour = 16'b11000_100111_01000; 
		6015: oled_colour = 16'b11001_101000_01001; 
		6016: oled_colour = 16'b11001_101000_01001; 
		6017: oled_colour = 16'b11000_100110_01000; 
		6018: oled_colour = 16'b11100_101111_01100; 
		6019: oled_colour = 16'b11011_101100_01011; 
		6020: oled_colour = 16'b11011_101100_01011; 
		6021: oled_colour = 16'b11010_101011_01010; 
		6022: oled_colour = 16'b11100_101110_01011; 
		6023: oled_colour = 16'b11001_101011_01010; 
		6024: oled_colour = 16'b11010_101010_01010; 
		6025: oled_colour = 16'b11011_101101_01011; 
		6026: oled_colour = 16'b11010_101001_01001; 
		6027: oled_colour = 16'b11100_101110_01011; 
		6028: oled_colour = 16'b11010_101001_01001; 
		6029: oled_colour = 16'b11000_100110_01000; 
		6030: oled_colour = 16'b11100_101110_01011; 
		6031: oled_colour = 16'b11011_101100_01011; 
		6032: oled_colour = 16'b11011_101101_01011; 
		6033: oled_colour = 16'b11010_101001_01001; 
		6034: oled_colour = 16'b11011_101100_01010; 
		6035: oled_colour = 16'b11011_101110_01011; 
		6036: oled_colour = 16'b11010_101011_01010; 
		6037: oled_colour = 16'b11011_101101_01011; 
		6038: oled_colour = 16'b11011_101100_01011; 
		6039: oled_colour = 16'b11100_101111_01100; 
		6040: oled_colour = 16'b11000_100110_01001; 
		6041: oled_colour = 16'b10111_100101_01000; 
		6042: oled_colour = 16'b11100_101111_01011; 
		6043: oled_colour = 16'b11011_101100_01010; 
		6044: oled_colour = 16'b11001_101001_01001; 
		6045: oled_colour = 16'b11011_101101_01011; 
		6046: oled_colour = 16'b11011_101110_01011; 
		6047: oled_colour = 16'b11001_101000_01001; 
		6048: oled_colour = 16'b10000_010111_00100; 
		6049: oled_colour = 16'b10000_010101_00011; 
		6050: oled_colour = 16'b10000_010101_00011; 
		6051: oled_colour = 16'b10000_010101_00011; 
		6052: oled_colour = 16'b10000_010101_00011; 
		6053: oled_colour = 16'b10000_010110_00011; 
		6054: oled_colour = 16'b10000_010101_00011; 
		6055: oled_colour = 16'b10000_010101_00011; 
		6056: oled_colour = 16'b10000_010101_00011; 
		6057: oled_colour = 16'b10000_010101_00011; 
		6058: oled_colour = 16'b10000_010101_00011; 
		6059: oled_colour = 16'b10000_010101_00011; 
		6060: oled_colour = 16'b10000_010110_00011; 
		6061: oled_colour = 16'b10000_010101_00011; 
		6062: oled_colour = 16'b10000_010101_00011; 
		6063: oled_colour = 16'b10000_010101_00011; 
		6064: oled_colour = 16'b10000_010101_00011; 
		6065: oled_colour = 16'b01111_010101_00011; 
		6066: oled_colour = 16'b10000_010101_00011; 
		6067: oled_colour = 16'b10000_010101_00011; 
		6068: oled_colour = 16'b10000_010101_00011; 
		6069: oled_colour = 16'b10000_010101_00011; 
		6070: oled_colour = 16'b10000_010110_00100; 
		6071: oled_colour = 16'b10001_010111_00100; 
		6072: oled_colour = 16'b10000_010101_00011; 
		6073: oled_colour = 16'b10000_010101_00011; 
		6074: oled_colour = 16'b10000_010101_00011; 
		6075: oled_colour = 16'b10000_010101_00011; 
		6076: oled_colour = 16'b10000_010101_00011; 
		6077: oled_colour = 16'b10000_010100_00011; 
		6078: oled_colour = 16'b10000_010101_00011; 
		6079: oled_colour = 16'b10000_010101_00011; 
		6080: oled_colour = 16'b10000_010101_00011; 
		6081: oled_colour = 16'b10000_010101_00011; 
		6082: oled_colour = 16'b01111_010101_00011; 
		6083: oled_colour = 16'b10000_010110_00100; 
		6084: oled_colour = 16'b10000_010101_00011; 
		6085: oled_colour = 16'b10000_010101_00011; 
		6086: oled_colour = 16'b10000_010101_00011; 
		6087: oled_colour = 16'b10000_010101_00011; 
		6088: oled_colour = 16'b10000_010101_00011; 
		6089: oled_colour = 16'b10000_010101_00011; 
		6090: oled_colour = 16'b10000_010101_00011; 
		6091: oled_colour = 16'b10000_010101_00011; 
		6092: oled_colour = 16'b10000_010101_00011; 
		6093: oled_colour = 16'b10000_010101_00011; 
		6094: oled_colour = 16'b01111_010100_00011; 
		6095: oled_colour = 16'b10000_010101_00011; 
		6096: oled_colour = 16'b10000_010101_00011; 
		6097: oled_colour = 16'b10000_010101_00011; 
		6098: oled_colour = 16'b10000_010101_00011; 
		6099: oled_colour = 16'b10000_010101_00011; 
		6100: oled_colour = 16'b10000_010101_00011; 
		6101: oled_colour = 16'b10000_010101_00011; 
		6102: oled_colour = 16'b10000_010101_00011; 
		6103: oled_colour = 16'b10000_010101_00011; 
		6104: oled_colour = 16'b10000_010101_00011; 
		6105: oled_colour = 16'b01111_010101_00011; 
		6106: oled_colour = 16'b10000_010101_00011; 
		6107: oled_colour = 16'b01111_010101_00011; 
		6108: oled_colour = 16'b01111_010100_00011; 
		6109: oled_colour = 16'b10000_010101_00011; 
		6110: oled_colour = 16'b10000_010110_00011; 
		6111: oled_colour = 16'b10000_010101_00011; 
		6112: oled_colour = 16'b10000_010101_00011; 
		6113: oled_colour = 16'b10000_010101_00011; 
		6114: oled_colour = 16'b10000_010101_00011; 
		6115: oled_colour = 16'b10000_010101_00011; 
		6116: oled_colour = 16'b10000_010101_00011; 
		6117: oled_colour = 16'b10000_010101_00011; 
		6118: oled_colour = 16'b10000_010110_00011; 
		6119: oled_colour = 16'b10000_010110_00011; 
		6120: oled_colour = 16'b10000_010100_00011; 
		6121: oled_colour = 16'b10000_010101_00011; 
		6122: oled_colour = 16'b10000_010101_00011; 
		6123: oled_colour = 16'b10000_010101_00011; 
		6124: oled_colour = 16'b10000_010101_00011; 
		6125: oled_colour = 16'b10000_010100_00011; 
		6126: oled_colour = 16'b10000_010101_00011; 
		6127: oled_colour = 16'b10000_010101_00011; 
		6128: oled_colour = 16'b10000_010101_00011; 
		6129: oled_colour = 16'b10000_010101_00011; 
		6130: oled_colour = 16'b10000_010101_00011; 
		6131: oled_colour = 16'b10001_010111_00100; 
		6132: oled_colour = 16'b10000_010101_00011; 
		6133: oled_colour = 16'b10000_010101_00011; 
		6134: oled_colour = 16'b10000_010101_00011; 
		6135: oled_colour = 16'b10000_010101_00011; 
		6136: oled_colour = 16'b10000_010101_00011; 
		6137: oled_colour = 16'b10000_010101_00011; 
		6138: oled_colour = 16'b10000_010101_00011; 
		6139: oled_colour = 16'b10000_010101_00011; 
		6140: oled_colour = 16'b01111_010101_00011; 
		6141: oled_colour = 16'b10000_010101_00011; 
		6142: oled_colour = 16'b10000_010110_00011; 
		6143: oled_colour = 16'b10000_010101_00011; 
		default: oled_colour = 16'b00000_000000_00000; 
	endcase
end

endmodule