module Gui_Inj2(
    input [12:0] pixel_index, 
    output reg [15:0] oled_colour 
); 

always@(pixel_index) 
begin
	case(pixel_index)
		2159: oled_colour = 16'b11111_111101_11111; 
		2160: oled_colour = 16'b11110_110110_11010; 
		2161: oled_colour = 16'b11100_110011_10100; 
		2162: oled_colour = 16'b11111_111100_11111; 
		2250: oled_colour = 16'b11100_110101_11011; 
		2251: oled_colour = 16'b11011_101111_10111; 
		2252: oled_colour = 16'b11101_110100_10111; 
		2253: oled_colour = 16'b11101_110011_10111; 
		2254: oled_colour = 16'b11001_101100_10100; 
		2255: oled_colour = 16'b10010_101001_10011; 
		2256: oled_colour = 16'b11010_101101_01100; 
		2257: oled_colour = 16'b11111_111000_00100; 
		2258: oled_colour = 16'b11101_110101_01010; 
		2259: oled_colour = 16'b11110_110111_10111; 
		2260: oled_colour = 16'b11111_111100_11111; 
		2344: oled_colour = 16'b11011_110001_11001; 
		2345: oled_colour = 16'b11011_101101_10100; 
		2346: oled_colour = 16'b11001_100100_10000; 
		2347: oled_colour = 16'b10111_100001_01110; 
		2348: oled_colour = 16'b11111_110101_10101; 
		2349: oled_colour = 16'b11110_110101_11001; 
		2350: oled_colour = 16'b11011_101011_10000; 
		2351: oled_colour = 16'b10010_110000_01111; 
		2352: oled_colour = 16'b11011_110010_01001; 
		2353: oled_colour = 16'b11111_110100_01010; 
		2354: oled_colour = 16'b11110_110110_00111; 
		2355: oled_colour = 16'b11110_110111_00100; 
		2356: oled_colour = 16'b11101_110100_01010; 
		2357: oled_colour = 16'b11110_110111_11010; 
		2358: oled_colour = 16'b11111_111110_11111; 
		2438: oled_colour = 16'b11011_110010_11001; 
		2439: oled_colour = 16'b11010_101011_10100; 
		2440: oled_colour = 16'b11011_101001_10000; 
		2441: oled_colour = 16'b11110_110110_11000; 
		2442: oled_colour = 16'b11110_101101_10001; 
		2443: oled_colour = 16'b11011_011110_01001; 
		2444: oled_colour = 16'b11100_100111_01111; 
		2445: oled_colour = 16'b11111_110110_10110; 
		2446: oled_colour = 16'b11100_101111_10100; 
		2447: oled_colour = 16'b10101_100101_01100; 
		2448: oled_colour = 16'b11101_110011_00110; 
		2449: oled_colour = 16'b11110_110110_01000; 
		2450: oled_colour = 16'b11110_110100_00111; 
		2451: oled_colour = 16'b11110_110011_01001; 
		2452: oled_colour = 16'b11110_110111_00110; 
		2453: oled_colour = 16'b11100_101110_01101; 
		2454: oled_colour = 16'b11011_101110_11001; 
		2455: oled_colour = 16'b11111_111110_11111; 
		2533: oled_colour = 16'b11011_110001_11000; 
		2534: oled_colour = 16'b11010_100100_01111; 
		2535: oled_colour = 16'b11101_101111_10100; 
		2536: oled_colour = 16'b11101_101101_10010; 
		2537: oled_colour = 16'b11110_110100_10100; 
		2538: oled_colour = 16'b11111_111001_11000; 
		2539: oled_colour = 16'b11011_100101_01110; 
		2540: oled_colour = 16'b11001_100001_01101; 
		2541: oled_colour = 16'b11110_101100_10000; 
		2542: oled_colour = 16'b11000_100111_01111; 
		2543: oled_colour = 16'b11000_100011_01101; 
		2544: oled_colour = 16'b11000_100101_01011; 
		2545: oled_colour = 16'b11011_101000_01100; 
		2546: oled_colour = 16'b11110_110010_01111; 
		2547: oled_colour = 16'b11101_110000_01010; 
		2548: oled_colour = 16'b11100_101100_01100; 
		2549: oled_colour = 16'b11101_101111_01000; 
		2550: oled_colour = 16'b11101_110011_10111; 
		2551: oled_colour = 16'b11111_111110_11111; 
		2629: oled_colour = 16'b11100_110011_11000; 
		2630: oled_colour = 16'b11101_101110_10010; 
		2631: oled_colour = 16'b11110_110011_10100; 
		2632: oled_colour = 16'b11011_100111_01111; 
		2633: oled_colour = 16'b11010_100110_01110; 
		2634: oled_colour = 16'b10100_100010_01011; 
		2635: oled_colour = 16'b01111_011001_00110; 
		2636: oled_colour = 16'b10000_010101_00101; 
		2637: oled_colour = 16'b10111_100110_01110; 
		2638: oled_colour = 16'b10111_101110_10001; 
		2639: oled_colour = 16'b11000_101010_10001; 
		2640: oled_colour = 16'b11001_100100_01110; 
		2641: oled_colour = 16'b11100_101110_10100; 
		2642: oled_colour = 16'b11011_101100_10100; 
		2643: oled_colour = 16'b11010_101001_10001; 
		2644: oled_colour = 16'b11001_101110_10100; 
		2645: oled_colour = 16'b11000_100001_01101; 
		2646: oled_colour = 16'b11011_101000_01110; 
		2647: oled_colour = 16'b11111_111110_11111; 
		2725: oled_colour = 16'b11100_110011_11001; 
		2726: oled_colour = 16'b11100_101010_01111; 
		2727: oled_colour = 16'b11110_110101_10100; 
		2728: oled_colour = 16'b11100_101000_10000; 
		2729: oled_colour = 16'b10001_010110_00110; 
		2730: oled_colour = 16'b00010_010001_00001; 
		2731: oled_colour = 16'b00010_010101_00001; 
		2732: oled_colour = 16'b00110_010101_00011; 
		2733: oled_colour = 16'b01001_011110_01001; 
		2734: oled_colour = 16'b10010_101010_10000; 
		2735: oled_colour = 16'b11001_101101_10000; 
		2736: oled_colour = 16'b11001_100011_01101; 
		2737: oled_colour = 16'b11101_101110_10011; 
		2738: oled_colour = 16'b11000_101000_10000; 
		2739: oled_colour = 16'b10010_100110_01101; 
		2740: oled_colour = 16'b11100_101011_10001; 
		2741: oled_colour = 16'b11101_110000_10101; 
		2742: oled_colour = 16'b11101_110001_10101; 
		2743: oled_colour = 16'b11000_100100_10000; 
		2744: oled_colour = 16'b11111_111101_11111; 
		2821: oled_colour = 16'b11110_111100_11111; 
		2822: oled_colour = 16'b11001_100111_10000; 
		2823: oled_colour = 16'b11111_111000_10111; 
		2824: oled_colour = 16'b11110_110000_10011; 
		2825: oled_colour = 16'b10101_011110_01010; 
		2826: oled_colour = 16'b01001_010110_00100; 
		2827: oled_colour = 16'b00111_010101_00010; 
		2828: oled_colour = 16'b01000_011011_00101; 
		2829: oled_colour = 16'b00110_010101_00010; 
		2830: oled_colour = 16'b01010_011100_01001; 
		2831: oled_colour = 16'b10101_101000_10001; 
		2832: oled_colour = 16'b10101_100110_01111; 
		2833: oled_colour = 16'b10110_100010_01110; 
		2834: oled_colour = 16'b10101_101011_10011; 
		2835: oled_colour = 16'b11001_110000_10111; 
		2836: oled_colour = 16'b11001_100010_01101; 
		2837: oled_colour = 16'b11110_110010_10011; 
		2838: oled_colour = 16'b11101_101111_10100; 
		2839: oled_colour = 16'b11011_101001_10000; 
		2840: oled_colour = 16'b11011_101110_10110; 
		2918: oled_colour = 16'b10000_100000_01100; 
		2919: oled_colour = 16'b11011_101100_10001; 
		2920: oled_colour = 16'b11111_111111_11101; 
		2921: oled_colour = 16'b11011_101011_10010; 
		2922: oled_colour = 16'b10000_100110_01110; 
		2923: oled_colour = 16'b01111_100111_01110; 
		2924: oled_colour = 16'b01111_100110_01110; 
		2925: oled_colour = 16'b01010_011100_00111; 
		2926: oled_colour = 16'b00101_010111_00100; 
		2927: oled_colour = 16'b10110_101111_10111; 
		2928: oled_colour = 16'b11110_111010_11101; 
		2929: oled_colour = 16'b11100_110111_11100; 
		2930: oled_colour = 16'b11111_111110_11111; 
		2932: oled_colour = 16'b11011_110010_11001; 
		2933: oled_colour = 16'b11001_100111_10001; 
		2934: oled_colour = 16'b11001_100010_01101; 
		2935: oled_colour = 16'b11101_101101_10010; 
		2936: oled_colour = 16'b11101_101111_10011; 
		2937: oled_colour = 16'b11011_101101_10110; 
		3014: oled_colour = 16'b10001_101001_10010; 
		3015: oled_colour = 16'b10100_100001_01100; 
		3016: oled_colour = 16'b11110_101111_10100; 
		3017: oled_colour = 16'b11100_101001_10001; 
		3018: oled_colour = 16'b11011_101011_10000; 
		3019: oled_colour = 16'b11001_101110_10001; 
		3020: oled_colour = 16'b01011_011110_01001; 
		3021: oled_colour = 16'b01000_011100_01000; 
		3022: oled_colour = 16'b01011_100001_01011; 
		3023: oled_colour = 16'b10000_100010_01011; 
		3024: oled_colour = 16'b11011_110011_11001; 
		3029: oled_colour = 16'b11011_110000_11000; 
		3030: oled_colour = 16'b11100_101111_10011; 
		3031: oled_colour = 16'b11111_111001_11000; 
		3032: oled_colour = 16'b11011_101001_10000; 
		3033: oled_colour = 16'b11010_101111_10111; 
		3110: oled_colour = 16'b11100_111001_11100; 
		3111: oled_colour = 16'b10110_100110_01111; 
		3112: oled_colour = 16'b11100_100100_01110; 
		3113: oled_colour = 16'b11110_101110_10001; 
		3114: oled_colour = 16'b11011_101100_10000; 
		3115: oled_colour = 16'b10001_100000_01010; 
		3116: oled_colour = 16'b01101_011011_00110; 
		3117: oled_colour = 16'b01001_011111_01001; 
		3118: oled_colour = 16'b10101_110110_10100; 
		3119: oled_colour = 16'b11001_110111_10110; 
		3120: oled_colour = 16'b01110_100100_01110; 
		3121: oled_colour = 16'b11100_111000_11100; 
		3124: oled_colour = 16'b11110_111010_11101; 
		3125: oled_colour = 16'b11011_101011_10100; 
		3126: oled_colour = 16'b11110_110101_10101; 
		3127: oled_colour = 16'b11101_110001_10011; 
		3128: oled_colour = 16'b11001_101001_10011; 
		3129: oled_colour = 16'b11111_111110_11111; 
		3206: oled_colour = 16'b11110_110111_11011; 
		3207: oled_colour = 16'b10101_011111_01011; 
		3208: oled_colour = 16'b11100_110001_10011; 
		3209: oled_colour = 16'b11110_110101_10110; 
		3210: oled_colour = 16'b11001_101001_01111; 
		3211: oled_colour = 16'b01100_100000_01100; 
		3212: oled_colour = 16'b01001_011100_01001; 
		3213: oled_colour = 16'b01011_100000_01010; 
		3214: oled_colour = 16'b11100_111111_11000; 
		3215: oled_colour = 16'b11101_111110_11010; 
		3216: oled_colour = 16'b11000_110111_10101; 
		3217: oled_colour = 16'b10011_101100_10011; 
		3218: oled_colour = 16'b11110_110111_11011; 
		3219: oled_colour = 16'b11010_100111_10010; 
		3220: oled_colour = 16'b11100_101101_10010; 
		3221: oled_colour = 16'b11101_110001_10010; 
		3222: oled_colour = 16'b11101_101110_10001; 
		3223: oled_colour = 16'b11001_101001_10010; 
		3224: oled_colour = 16'b11111_111101_11111; 
		3302: oled_colour = 16'b11001_110001_11000; 
		3303: oled_colour = 16'b01001_011111_01000; 
		3304: oled_colour = 16'b10111_101110_10001; 
		3305: oled_colour = 16'b11001_100110_01110; 
		3306: oled_colour = 16'b11001_101001_01110; 
		3307: oled_colour = 16'b10011_100110_01111; 
		3308: oled_colour = 16'b11100_111010_11110; 
		3309: oled_colour = 16'b01111_100100_01110; 
		3310: oled_colour = 16'b01110_101001_01110; 
		3311: oled_colour = 16'b10100_110110_10011; 
		3312: oled_colour = 16'b11110_111111_11010; 
		3313: oled_colour = 16'b10100_110011_10010; 
		3314: oled_colour = 16'b10101_101010_10100; 
		3315: oled_colour = 16'b11100_110000_10111; 
		3316: oled_colour = 16'b11100_101110_10011; 
		3317: oled_colour = 16'b11111_111101_11010; 
		3318: oled_colour = 16'b11011_101001_01111; 
		3319: oled_colour = 16'b11110_111001_11101; 
		3398: oled_colour = 16'b11110_111101_11110; 
		3399: oled_colour = 16'b01101_100011_01101; 
		3400: oled_colour = 16'b01011_100001_01011; 
		3401: oled_colour = 16'b11000_110110_10011; 
		3402: oled_colour = 16'b11011_110100_10010; 
		3403: oled_colour = 16'b10011_100110_01111; 
		3404: oled_colour = 16'b11110_111101_11111; 
		3406: oled_colour = 16'b01110_100001_01101; 
		3407: oled_colour = 16'b10001_100111_01101; 
		3408: oled_colour = 16'b11000_111001_10101; 
		3409: oled_colour = 16'b10010_101010_01110; 
		3410: oled_colour = 16'b10101_101001_10011; 
		3411: oled_colour = 16'b11100_101101_10101; 
		3412: oled_colour = 16'b11010_100110_01111; 
		3413: oled_colour = 16'b11011_101011_10010; 
		3414: oled_colour = 16'b11011_101110_10110; 
		3496: oled_colour = 16'b01011_100001_01100; 
		3497: oled_colour = 16'b10011_110101_10010; 
		3498: oled_colour = 16'b10111_111001_10100; 
		3499: oled_colour = 16'b10100_100011_01110; 
		3500: oled_colour = 16'b11111_111011_11110; 
		3502: oled_colour = 16'b10111_101010_10011; 
		3503: oled_colour = 16'b10110_011100_01010; 
		3504: oled_colour = 16'b11011_101001_10000; 
		3505: oled_colour = 16'b10001_011010_01000; 
		3506: oled_colour = 16'b10000_011111_01100; 
		3507: oled_colour = 16'b11101_110111_11100; 
		3508: oled_colour = 16'b11100_110011_11001; 
		3509: oled_colour = 16'b11101_110101_11010; 
		3591: oled_colour = 16'b11110_111100_11110; 
		3592: oled_colour = 16'b01110_011010_01000; 
		3593: oled_colour = 16'b01110_100100_01101; 
		3594: oled_colour = 16'b01010_100011_01100; 
		3595: oled_colour = 16'b01000_011010_00110; 
		3596: oled_colour = 16'b11110_111100_11110; 
		3598: oled_colour = 16'b11000_110010_10111; 
		3599: oled_colour = 16'b01000_010110_00100; 
		3600: oled_colour = 16'b10001_100101_01110; 
		3601: oled_colour = 16'b01111_100111_01111; 
		3602: oled_colour = 16'b01010_011110_01010; 
		3603: oled_colour = 16'b11111_111110_11111; 
		3687: oled_colour = 16'b11001_110000_10111; 
		3688: oled_colour = 16'b01101_010111_00111; 
		3689: oled_colour = 16'b10001_011101_01010; 
		3690: oled_colour = 16'b00110_011001_00101; 
		3691: oled_colour = 16'b01000_011010_00110; 
		3692: oled_colour = 16'b11110_111100_11110; 
		3694: oled_colour = 16'b11101_111010_11101; 
		3695: oled_colour = 16'b00111_010011_00010; 
		3696: oled_colour = 16'b01001_011101_01001; 
		3697: oled_colour = 16'b01110_100010_01101; 
		3698: oled_colour = 16'b01011_010111_00110; 
		3699: oled_colour = 16'b11101_111010_11101; 
		3783: oled_colour = 16'b11000_110000_10110; 
		3784: oled_colour = 16'b01000_011001_00110; 
		3785: oled_colour = 16'b01101_100010_01101; 
		3786: oled_colour = 16'b01101_011100_01001; 
		3787: oled_colour = 16'b10011_100001_01110; 
		3791: oled_colour = 16'b01101_011101_01001; 
		3792: oled_colour = 16'b01001_011001_00101; 
		3793: oled_colour = 16'b01000_010111_00100; 
		3794: oled_colour = 16'b01111_100100_01110; 
		3879: oled_colour = 16'b11101_111010_11101; 
		3880: oled_colour = 16'b01100_011011_00111; 
		3881: oled_colour = 16'b01100_100000_01011; 
		3882: oled_colour = 16'b01010_011001_00110; 
		3883: oled_colour = 16'b11010_110100_11001; 
		3887: oled_colour = 16'b10111_101000_10011; 
		3888: oled_colour = 16'b10101_011010_01000; 
		3889: oled_colour = 16'b10110_100000_01100; 
		3890: oled_colour = 16'b11111_111110_11111; 
		3975: oled_colour = 16'b11111_111110_11111; 
		3976: oled_colour = 16'b10101_100000_01100; 
		3977: oled_colour = 16'b10011_011010_00111; 
		3978: oled_colour = 16'b11001_110001_11000; 
		3982: oled_colour = 16'b11111_111110_11111; 
		3983: oled_colour = 16'b10001_011010_01001; 
		3984: oled_colour = 16'b01101_001111_00001; 
		3985: oled_colour = 16'b10011_011101_01011; 
		3986: oled_colour = 16'b11100_110111_11100; 
		3987: oled_colour = 16'b11111_111110_11111; 
		4071: oled_colour = 16'b11100_110111_11011; 
		4072: oled_colour = 16'b10011_011100_01001; 
		4073: oled_colour = 16'b10011_011011_00111; 
		4074: oled_colour = 16'b11000_101101_10101; 
		4079: oled_colour = 16'b11000_101010_10011; 
		4080: oled_colour = 16'b01111_010111_00110; 
		4081: oled_colour = 16'b10000_010101_00100; 
		4082: oled_colour = 16'b11000_100001_01101; 
		4083: oled_colour = 16'b10101_011111_01101; 
		4084: oled_colour = 16'b11101_111000_11100; 
		4167: oled_colour = 16'b11001_101110_10110; 
		4168: oled_colour = 16'b10101_011100_01001; 
		4169: oled_colour = 16'b10100_011011_01001; 
		4170: oled_colour = 16'b10110_100111_10001; 
		4176: oled_colour = 16'b11111_111101_11111; 
		4177: oled_colour = 16'b11011_101100_10100; 
		4178: oled_colour = 16'b11110_101110_10010; 
		4179: oled_colour = 16'b11000_100011_01111; 
		4180: oled_colour = 16'b11101_110110_11011; 
		4263: oled_colour = 16'b11000_100111_10010; 
		4264: oled_colour = 16'b11010_100011_01100; 
		4265: oled_colour = 16'b11000_011111_01011; 
		4266: oled_colour = 16'b10101_100000_01110; 
		4274: oled_colour = 16'b11111_111110_11111; 
		4359: oled_colour = 16'b11110_111001_11100; 
		4360: oled_colour = 16'b11101_110100_11001; 
		4361: oled_colour = 16'b11101_110101_11001; 
		4362: oled_colour = 16'b11101_110111_11011; 
		default: oled_colour = 16'b00000_000000_00000; 
	endcase
end

endmodule