module Gui_Punch3(
    input [12:0] pixel_index, 
    output reg [15:0] oled_colour 
); 

always@(pixel_index) 
begin
	case(pixel_index)
		1773: oled_colour = 16'b11111_111110_11111; 
		1868: oled_colour = 16'b11111_111101_11111; 
		1869: oled_colour = 16'b11101_110011_11001; 
		1870: oled_colour = 16'b11100_101111_10000; 
		1871: oled_colour = 16'b11101_110100_01111; 
		1872: oled_colour = 16'b11110_110111_01100; 
		1873: oled_colour = 16'b11110_111001_01000; 
		1874: oled_colour = 16'b11110_110110_01011; 
		1875: oled_colour = 16'b11110_110111_01011; 
		1876: oled_colour = 16'b11101_110001_10000; 
		1877: oled_colour = 16'b11110_111001_11101; 
		1966: oled_colour = 16'b11101_110111_11010; 
		1967: oled_colour = 16'b11100_101100_01001; 
		1968: oled_colour = 16'b11101_110001_01010; 
		1969: oled_colour = 16'b11011_101101_01010; 
		1970: oled_colour = 16'b11110_110001_01010; 
		1971: oled_colour = 16'b11101_110001_01001; 
		1972: oled_colour = 16'b11110_111000_11010; 
		2058: oled_colour = 16'b11111_111100_11111; 
		2059: oled_colour = 16'b11110_110110_11010; 
		2060: oled_colour = 16'b11000_101001_10001; 
		2061: oled_colour = 16'b10010_101011_10010; 
		2062: oled_colour = 16'b11000_101000_10000; 
		2063: oled_colour = 16'b11010_101000_01111; 
		2064: oled_colour = 16'b11011_101001_10000; 
		2065: oled_colour = 16'b11011_101011_10010; 
		2066: oled_colour = 16'b11011_110000_10110; 
		2067: oled_colour = 16'b11100_110000_10111; 
		2153: oled_colour = 16'b11110_110111_11011; 
		2154: oled_colour = 16'b11101_110011_10110; 
		2155: oled_colour = 16'b11110_111000_11000; 
		2156: oled_colour = 16'b11110_110000_10010; 
		2157: oled_colour = 16'b10011_100111_01110; 
		2158: oled_colour = 16'b10011_011111_01010; 
		2159: oled_colour = 16'b10011_011100_01010; 
		2160: oled_colour = 16'b11001_100100_01110; 
		2161: oled_colour = 16'b11101_101101_10010; 
		2162: oled_colour = 16'b11001_101011_10010; 
		2163: oled_colour = 16'b11011_101100_10010; 
		2164: oled_colour = 16'b11110_111000_11011; 
		2165: oled_colour = 16'b11111_111110_11111; 
		2249: oled_colour = 16'b11100_110010_11000; 
		2250: oled_colour = 16'b11010_011110_01000; 
		2251: oled_colour = 16'b10111_100100_10001; 
		2252: oled_colour = 16'b11011_101000_10000; 
		2253: oled_colour = 16'b11000_100000_01100; 
		2254: oled_colour = 16'b11011_101100_10010; 
		2255: oled_colour = 16'b10110_100011_01100; 
		2256: oled_colour = 16'b10001_010110_00110; 
		2257: oled_colour = 16'b11001_100100_01101; 
		2258: oled_colour = 16'b11000_100110_01101; 
		2259: oled_colour = 16'b10101_100001_01100; 
		2260: oled_colour = 16'b11100_100111_01111; 
		2261: oled_colour = 16'b11011_101001_10011; 
		2264: oled_colour = 16'b11110_111011_11110; 
		2265: oled_colour = 16'b11011_101110_10110; 
		2266: oled_colour = 16'b11101_110001_10110; 
		2267: oled_colour = 16'b11100_101110_10101; 
		2268: oled_colour = 16'b11011_101101_10101; 
		2345: oled_colour = 16'b11010_101100_10100; 
		2346: oled_colour = 16'b11011_100110_01110; 
		2347: oled_colour = 16'b11110_101111_10010; 
		2348: oled_colour = 16'b11000_100010_01101; 
		2349: oled_colour = 16'b11000_100000_01100; 
		2350: oled_colour = 16'b11111_110010_10100; 
		2351: oled_colour = 16'b11011_101011_10001; 
		2352: oled_colour = 16'b10110_011110_01010; 
		2353: oled_colour = 16'b10010_011001_01000; 
		2354: oled_colour = 16'b10001_011101_01001; 
		2355: oled_colour = 16'b10001_011101_01010; 
		2356: oled_colour = 16'b11011_101000_10000; 
		2357: oled_colour = 16'b11011_101100_10010; 
		2358: oled_colour = 16'b11010_101111_10111; 
		2359: oled_colour = 16'b11011_110010_11001; 
		2360: oled_colour = 16'b11011_101001_10000; 
		2361: oled_colour = 16'b11101_101010_01111; 
		2362: oled_colour = 16'b11011_101011_01111; 
		2363: oled_colour = 16'b11000_011111_01011; 
		2364: oled_colour = 16'b11001_100111_10001; 
		2441: oled_colour = 16'b11011_101101_10100; 
		2442: oled_colour = 16'b11110_110010_10100; 
		2443: oled_colour = 16'b11100_101100_10001; 
		2444: oled_colour = 16'b11010_100100_01110; 
		2445: oled_colour = 16'b11101_101010_10000; 
		2446: oled_colour = 16'b10111_100001_01100; 
		2447: oled_colour = 16'b10000_100010_01101; 
		2448: oled_colour = 16'b10010_101010_10000; 
		2449: oled_colour = 16'b01111_100101_01101; 
		2450: oled_colour = 16'b01011_100011_01011; 
		2451: oled_colour = 16'b10010_100001_01100; 
		2452: oled_colour = 16'b11111_110000_10001; 
		2453: oled_colour = 16'b11101_101110_10010; 
		2454: oled_colour = 16'b11000_100010_01101; 
		2455: oled_colour = 16'b11010_100110_01111; 
		2456: oled_colour = 16'b11101_101101_10001; 
		2457: oled_colour = 16'b11010_101100_10100; 
		2458: oled_colour = 16'b11101_110100_11001; 
		2459: oled_colour = 16'b11101_110011_11001; 
		2460: oled_colour = 16'b11111_111110_11111; 
		2537: oled_colour = 16'b11101_110011_11000; 
		2538: oled_colour = 16'b11101_101111_10001; 
		2539: oled_colour = 16'b11100_101110_10010; 
		2540: oled_colour = 16'b11110_110001_10011; 
		2541: oled_colour = 16'b11011_101001_01111; 
		2542: oled_colour = 16'b01001_011000_00110; 
		2543: oled_colour = 16'b00110_011011_00110; 
		2544: oled_colour = 16'b00100_010111_00011; 
		2545: oled_colour = 16'b01000_011011_01000; 
		2546: oled_colour = 16'b10001_101001_10010; 
		2547: oled_colour = 16'b11011_110100_11010; 
		2548: oled_colour = 16'b11011_101100_10101; 
		2549: oled_colour = 16'b11011_100101_01111; 
		2550: oled_colour = 16'b11101_101011_01111; 
		2551: oled_colour = 16'b11111_110011_10100; 
		2552: oled_colour = 16'b11011_101010_10010; 
		2553: oled_colour = 16'b11110_111011_11110; 
		2633: oled_colour = 16'b11101_110110_11011; 
		2634: oled_colour = 16'b11100_101101_10001; 
		2635: oled_colour = 16'b11111_111001_11001; 
		2636: oled_colour = 16'b11111_110101_10111; 
		2637: oled_colour = 16'b10000_011011_01000; 
		2638: oled_colour = 16'b00010_010100_00001; 
		2639: oled_colour = 16'b00010_010011_00001; 
		2640: oled_colour = 16'b00110_011000_00101; 
		2641: oled_colour = 16'b11001_110101_11010; 
		2645: oled_colour = 16'b11110_111001_11101; 
		2646: oled_colour = 16'b11100_101111_10110; 
		2647: oled_colour = 16'b11101_110001_10110; 
		2648: oled_colour = 16'b11101_110110_11011; 
		2729: oled_colour = 16'b11110_111100_11110; 
		2730: oled_colour = 16'b10100_100000_01100; 
		2731: oled_colour = 16'b11010_101000_01111; 
		2732: oled_colour = 16'b10011_011001_00111; 
		2733: oled_colour = 16'b01100_010010_00011; 
		2734: oled_colour = 16'b10000_011111_01011; 
		2735: oled_colour = 16'b01111_011110_01001; 
		2736: oled_colour = 16'b10010_100101_01111; 
		2825: oled_colour = 16'b11100_111000_11100; 
		2826: oled_colour = 16'b01111_011110_01010; 
		2827: oled_colour = 16'b10010_101010_01110; 
		2828: oled_colour = 16'b01100_011100_00110; 
		2829: oled_colour = 16'b01110_010111_00110; 
		2830: oled_colour = 16'b01101_100101_01100; 
		2831: oled_colour = 16'b01110_011110_01000; 
		2832: oled_colour = 16'b01110_011100_01010; 
		2833: oled_colour = 16'b11110_111101_11111; 
		2920: oled_colour = 16'b11111_111110_11111; 
		2921: oled_colour = 16'b11001_110100_11001; 
		2922: oled_colour = 16'b01111_011101_01001; 
		2923: oled_colour = 16'b10101_101010_01110; 
		2924: oled_colour = 16'b11000_101111_01111; 
		2925: oled_colour = 16'b10110_100101_01100; 
		2926: oled_colour = 16'b01010_100100_01010; 
		2927: oled_colour = 16'b01101_100001_01001; 
		2928: oled_colour = 16'b10001_011100_01010; 
		2929: oled_colour = 16'b11100_111001_11101; 
		3016: oled_colour = 16'b11100_111010_11100; 
		3017: oled_colour = 16'b10110_110010_10101; 
		3018: oled_colour = 16'b10000_101101_10010; 
		3019: oled_colour = 16'b10110_111010_10100; 
		3020: oled_colour = 16'b11100_111011_11000; 
		3021: oled_colour = 16'b10101_101111_10010; 
		3022: oled_colour = 16'b00111_011100_00110; 
		3023: oled_colour = 16'b01111_100111_01100; 
		3024: oled_colour = 16'b10000_100101_01101; 
		3025: oled_colour = 16'b10011_100101_01111; 
		3026: oled_colour = 16'b11110_111010_11101; 
		3112: oled_colour = 16'b11100_111010_11100; 
		3113: oled_colour = 16'b10110_110100_10110; 
		3114: oled_colour = 16'b10101_101001_10001; 
		3115: oled_colour = 16'b11101_110010_10011; 
		3116: oled_colour = 16'b11111_111000_11000; 
		3117: oled_colour = 16'b11010_111000_10110; 
		3118: oled_colour = 16'b00110_011011_00101; 
		3119: oled_colour = 16'b01010_010101_00100; 
		3120: oled_colour = 16'b11001_101001_10001; 
		3121: oled_colour = 16'b11110_110011_10110; 
		3122: oled_colour = 16'b11100_101110_10100; 
		3123: oled_colour = 16'b11101_110101_11010; 
		3208: oled_colour = 16'b11110_111000_11100; 
		3209: oled_colour = 16'b11101_110001_10100; 
		3210: oled_colour = 16'b11100_101100_10011; 
		3211: oled_colour = 16'b11110_110010_10101; 
		3212: oled_colour = 16'b11111_111001_11000; 
		3213: oled_colour = 16'b11001_111000_10110; 
		3214: oled_colour = 16'b01010_011100_01000; 
		3215: oled_colour = 16'b01001_010100_00100; 
		3216: oled_colour = 16'b10110_110001_10011; 
		3217: oled_colour = 16'b11110_110111_10100; 
		3218: oled_colour = 16'b11100_110111_10011; 
		3219: oled_colour = 16'b11010_100111_01111; 
		3220: oled_colour = 16'b11011_110101_11011; 
		3304: oled_colour = 16'b11110_111000_11100; 
		3305: oled_colour = 16'b11100_110100_11000; 
		3306: oled_colour = 16'b11011_101100_10011; 
		3307: oled_colour = 16'b11101_101110_10000; 
		3308: oled_colour = 16'b11111_111011_11011; 
		3309: oled_colour = 16'b10111_110110_10100; 
		3310: oled_colour = 16'b11001_110101_11001; 
		3311: oled_colour = 16'b10010_101000_10001; 
		3312: oled_colour = 16'b10101_101101_10011; 
		3313: oled_colour = 16'b11001_111010_10111; 
		3314: oled_colour = 16'b11100_110100_10010; 
		3315: oled_colour = 16'b11101_111001_10100; 
		3316: oled_colour = 16'b10110_110101_10011; 
		3317: oled_colour = 16'b11101_111011_11110; 
		3401: oled_colour = 16'b10100_110000_10110; 
		3402: oled_colour = 16'b10000_101001_01111; 
		3403: oled_colour = 16'b11010_111001_10110; 
		3404: oled_colour = 16'b11111_111010_10111; 
		3405: oled_colour = 16'b10111_110010_10011; 
		3406: oled_colour = 16'b11011_111001_11100; 
		3408: oled_colour = 16'b10000_100100_01111; 
		3409: oled_colour = 16'b00111_011011_00111; 
		3410: oled_colour = 16'b10001_101110_10000; 
		3411: oled_colour = 16'b11001_111100_10101; 
		3412: oled_colour = 16'b10111_110001_10000; 
		3413: oled_colour = 16'b11100_110111_11011; 
		3496: oled_colour = 16'b11110_110110_11010; 
		3497: oled_colour = 16'b01110_010110_00101; 
		3498: oled_colour = 16'b01010_011000_00110; 
		3499: oled_colour = 16'b10011_101100_10000; 
		3500: oled_colour = 16'b11010_111100_10101; 
		3501: oled_colour = 16'b10100_110010_10100; 
		3503: oled_colour = 16'b11011_110100_11001; 
		3504: oled_colour = 16'b01110_010101_00101; 
		3505: oled_colour = 16'b10001_100111_01111; 
		3506: oled_colour = 16'b10110_111000_10100; 
		3507: oled_colour = 16'b11010_111000_10011; 
		3508: oled_colour = 16'b10011_100011_01101; 
		3509: oled_colour = 16'b11101_111010_11101; 
		3591: oled_colour = 16'b11111_111101_11111; 
		3592: oled_colour = 16'b10111_101001_10010; 
		3593: oled_colour = 16'b11001_100011_01101; 
		3594: oled_colour = 16'b10111_101111_10000; 
		3595: oled_colour = 16'b11010_111000_10100; 
		3596: oled_colour = 16'b10011_101110_01111; 
		3597: oled_colour = 16'b10101_101111_10110; 
		3599: oled_colour = 16'b10101_101110_10101; 
		3600: oled_colour = 16'b01011_010110_00101; 
		3601: oled_colour = 16'b11010_101001_10001; 
		3602: oled_colour = 16'b11111_110110_10110; 
		3603: oled_colour = 16'b11011_101110_10010; 
		3604: oled_colour = 16'b11011_110000_11000; 
		3687: oled_colour = 16'b11011_110011_11000; 
		3688: oled_colour = 16'b01100_011001_00111; 
		3689: oled_colour = 16'b11010_110010_11000; 
		3690: oled_colour = 16'b11110_110101_10101; 
		3691: oled_colour = 16'b11000_101001_01110; 
		3692: oled_colour = 16'b10011_100000_01101; 
		3693: oled_colour = 16'b11111_111011_11110; 
		3695: oled_colour = 16'b11011_111000_11100; 
		3696: oled_colour = 16'b00101_010111_00100; 
		3697: oled_colour = 16'b01010_011101_01000; 
		3698: oled_colour = 16'b01110_011100_01000; 
		3699: oled_colour = 16'b10010_100110_10000; 
		3783: oled_colour = 16'b11010_101110_10101; 
		3784: oled_colour = 16'b01011_010100_00011; 
		3785: oled_colour = 16'b01001_011101_01001; 
		3786: oled_colour = 16'b01101_100011_01101; 
		3787: oled_colour = 16'b10000_100011_01111; 
		3788: oled_colour = 16'b11101_111001_11101; 
		3791: oled_colour = 16'b11111_111100_11111; 
		3792: oled_colour = 16'b10101_011111_01100; 
		3793: oled_colour = 16'b10111_100001_01011; 
		3794: oled_colour = 16'b01101_010101_00101; 
		3795: oled_colour = 16'b11001_110010_11000; 
		3879: oled_colour = 16'b10010_011110_01011; 
		3880: oled_colour = 16'b10011_011010_00111; 
		3881: oled_colour = 16'b10001_011010_00111; 
		3882: oled_colour = 16'b10111_101100_10100; 
		3888: oled_colour = 16'b10001_011100_01010; 
		3889: oled_colour = 16'b01110_010001_00010; 
		3890: oled_colour = 16'b10100_011100_01010; 
		3891: oled_colour = 16'b11111_111110_11111; 
		3974: oled_colour = 16'b11001_110000_10111; 
		3975: oled_colour = 16'b01110_010011_00011; 
		3976: oled_colour = 16'b10001_011001_00110; 
		3977: oled_colour = 16'b10100_100011_01111; 
		3984: oled_colour = 16'b10101_100000_01110; 
		3985: oled_colour = 16'b01101_010010_00010; 
		3986: oled_colour = 16'b10000_010111_00110; 
		3987: oled_colour = 16'b11010_110000_10111; 
		4070: oled_colour = 16'b10011_011110_01100; 
		4071: oled_colour = 16'b11010_100110_01111; 
		4072: oled_colour = 16'b10100_011100_01001; 
		4073: oled_colour = 16'b11001_110000_10111; 
		4079: oled_colour = 16'b11110_111100_11110; 
		4080: oled_colour = 16'b10111_011111_01101; 
		4081: oled_colour = 16'b10010_011000_00110; 
		4082: oled_colour = 16'b01011_001101_00001; 
		4083: oled_colour = 16'b10001_010101_00110; 
		4084: oled_colour = 16'b11001_100110_10001; 
		4085: oled_colour = 16'b11101_110110_11011; 
		4165: oled_colour = 16'b11111_111101_11111; 
		4166: oled_colour = 16'b10110_100000_01101; 
		4167: oled_colour = 16'b11001_100101_01111; 
		4168: oled_colour = 16'b10101_011110_01100; 
		4169: oled_colour = 16'b11101_111000_11100; 
		4176: oled_colour = 16'b11100_110100_11000; 
		4177: oled_colour = 16'b11011_110001_10111; 
		4178: oled_colour = 16'b11000_101100_10100; 
		4179: oled_colour = 16'b10111_100011_01111; 
		4180: oled_colour = 16'b11010_101000_10001; 
		4181: oled_colour = 16'b11010_101001_10010; 
		4182: oled_colour = 16'b11101_111000_11100; 
		4262: oled_colour = 16'b11111_111100_11111; 
		4263: oled_colour = 16'b11100_110101_11001; 
		4264: oled_colour = 16'b11101_110111_11011; 
		4276: oled_colour = 16'b11111_111110_11111; 
		4277: oled_colour = 16'b11111_111110_11111; 
		default: oled_colour = 16'b00000_000000_00000; 
	endcase
end

endmodule