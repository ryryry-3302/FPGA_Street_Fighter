module Gui_Sp3(
    input [12:0] pixel_index, 
    output reg [15:0] oled_colour 
); 

always@(pixel_index) 
begin
	case(pixel_index)
		1968: oled_colour = 16'b11010_101001_01011; 
		1969: oled_colour = 16'b11111_111000_01001; 
		1970: oled_colour = 16'b11111_111010_00101; 
		1971: oled_colour = 16'b11111_111100_01001; 
		1972: oled_colour = 16'b11111_111011_01111; 
		1973: oled_colour = 16'b11110_110001_01100; 
		2061: oled_colour = 16'b01000_011011_00111; 
		2062: oled_colour = 16'b01110_011110_01000; 
		2063: oled_colour = 16'b10110_100001_01100; 
		2064: oled_colour = 16'b11010_101010_01011; 
		2065: oled_colour = 16'b11111_111010_00101; 
		2066: oled_colour = 16'b11101_110111_00100; 
		2067: oled_colour = 16'b11110_110100_01001; 
		2068: oled_colour = 16'b11111_110111_01011; 
		2069: oled_colour = 16'b11111_110011_01011; 
		2070: oled_colour = 16'b11011_101011_01010; 
		2155: oled_colour = 16'b01000_011010_00111; 
		2156: oled_colour = 16'b01100_100100_01100; 
		2157: oled_colour = 16'b01100_100101_01110; 
		2158: oled_colour = 16'b01111_100010_01011; 
		2159: oled_colour = 16'b10100_100001_01010; 
		2160: oled_colour = 16'b11000_100101_01011; 
		2161: oled_colour = 16'b11011_101111_01010; 
		2162: oled_colour = 16'b11100_101011_01011; 
		2163: oled_colour = 16'b11001_100101_10000; 
		2164: oled_colour = 16'b11010_101101_10011; 
		2165: oled_colour = 16'b11100_101100_10000; 
		2166: oled_colour = 16'b11101_101010_10000; 
		2167: oled_colour = 16'b11111_110011_10011; 
		2168: oled_colour = 16'b11101_110001_10010; 
		2169: oled_colour = 16'b11100_101110_10001; 
		2251: oled_colour = 16'b01111_101011_10000; 
		2252: oled_colour = 16'b01111_101100_10000; 
		2253: oled_colour = 16'b10100_101101_10010; 
		2254: oled_colour = 16'b11001_101010_10000; 
		2255: oled_colour = 16'b11010_101110_10010; 
		2256: oled_colour = 16'b11011_101100_10011; 
		2257: oled_colour = 16'b11000_100101_01101; 
		2258: oled_colour = 16'b11001_100010_01101; 
		2259: oled_colour = 16'b11011_101110_10011; 
		2260: oled_colour = 16'b11001_101001_10001; 
		2261: oled_colour = 16'b10111_100011_01101; 
		2262: oled_colour = 16'b11001_100011_01101; 
		2263: oled_colour = 16'b11111_110010_10100; 
		2264: oled_colour = 16'b11111_110111_10110; 
		2265: oled_colour = 16'b11111_110111_10101; 
		2266: oled_colour = 16'b11111_111001_11000; 
		2267: oled_colour = 16'b11100_101101_10010; 
		2346: oled_colour = 16'b01001_011101_01000; 
		2347: oled_colour = 16'b01100_100010_01100; 
		2348: oled_colour = 16'b10001_101001_01111; 
		2349: oled_colour = 16'b11101_101110_10011; 
		2350: oled_colour = 16'b11110_101111_10001; 
		2351: oled_colour = 16'b11111_111011_11001; 
		2352: oled_colour = 16'b11101_111100_11111; 
		2353: oled_colour = 16'b11010_100110_01110; 
		2354: oled_colour = 16'b10001_010110_00111; 
		2355: oled_colour = 16'b11100_101001_01111; 
		2356: oled_colour = 16'b11011_101110_10001; 
		2360: oled_colour = 16'b11001_100101_01110; 
		2361: oled_colour = 16'b11010_100110_01110; 
		2362: oled_colour = 16'b11011_101010_10000; 
		2363: oled_colour = 16'b11101_101011_10001; 
		2364: oled_colour = 16'b11111_101110_10001; 
		2365: oled_colour = 16'b11111_110001_10010; 
		2366: oled_colour = 16'b11100_101100_10000; 
		2442: oled_colour = 16'b00101_011000_00011; 
		2443: oled_colour = 16'b00101_010111_00100; 
		2444: oled_colour = 16'b10110_100101_01101; 
		2445: oled_colour = 16'b11111_110011_10101; 
		2446: oled_colour = 16'b11100_101001_10000; 
		2447: oled_colour = 16'b11011_100101_01101; 
		2448: oled_colour = 16'b10110_011000_01010; 
		2449: oled_colour = 16'b11001_011101_01010; 
		2450: oled_colour = 16'b11000_100101_01101; 
		2459: oled_colour = 16'b11010_100110_01110; 
		2460: oled_colour = 16'b11010_100100_01110; 
		2461: oled_colour = 16'b11001_101000_01110; 
		2462: oled_colour = 16'b11000_100011_01101; 
		2537: oled_colour = 16'b00011_010101_00001; 
		2538: oled_colour = 16'b00011_010101_00001; 
		2539: oled_colour = 16'b00010_010100_00001; 
		2540: oled_colour = 16'b10011_011011_01001; 
		2541: oled_colour = 16'b11000_011111_01100; 
		2542: oled_colour = 16'b10110_011101_01011; 
		2543: oled_colour = 16'b11011_100001_01100; 
		2544: oled_colour = 16'b11101_101000_01111; 
		2545: oled_colour = 16'b11100_101110_10100; 
		2546: oled_colour = 16'b11111_110010_10100; 
		2547: oled_colour = 16'b11111_110110_10110; 
		2556: oled_colour = 16'b11011_100111_01111; 
		2557: oled_colour = 16'b10111_100001_01100; 
		2633: oled_colour = 16'b00011_010100_00001; 
		2634: oled_colour = 16'b00011_010101_00001; 
		2635: oled_colour = 16'b00011_010101_00010; 
		2636: oled_colour = 16'b01011_011000_00110; 
		2637: oled_colour = 16'b10100_011011_01010; 
		2638: oled_colour = 16'b10000_011000_00111; 
		2639: oled_colour = 16'b10110_100001_01100; 
		2640: oled_colour = 16'b11111_110011_10100; 
		2641: oled_colour = 16'b11111_111001_11001; 
		2642: oled_colour = 16'b11110_110100_10110; 
		2643: oled_colour = 16'b11110_110011_10011; 
		2644: oled_colour = 16'b11100_101010_10000; 
		2651: oled_colour = 16'b11010_100101_01110; 
		2652: oled_colour = 16'b11110_110000_10010; 
		2653: oled_colour = 16'b11111_110011_10011; 
		2654: oled_colour = 16'b11100_101010_10000; 
		2729: oled_colour = 16'b00100_010110_00001; 
		2730: oled_colour = 16'b00010_010100_00001; 
		2731: oled_colour = 16'b00011_010100_00001; 
		2732: oled_colour = 16'b00100_010111_00010; 
		2733: oled_colour = 16'b01000_011001_00101; 
		2734: oled_colour = 16'b01000_011010_00111; 
		2737: oled_colour = 16'b11010_100100_01101; 
		2738: oled_colour = 16'b11111_110000_10011; 
		2739: oled_colour = 16'b11110_110000_10010; 
		2740: oled_colour = 16'b11100_101011_01111; 
		2741: oled_colour = 16'b11110_110000_10100; 
		2742: oled_colour = 16'b11111_110011_10101; 
		2743: oled_colour = 16'b11111_110100_10101; 
		2744: oled_colour = 16'b11111_110101_10100; 
		2745: oled_colour = 16'b11111_110011_10010; 
		2746: oled_colour = 16'b11111_110000_10010; 
		2747: oled_colour = 16'b11111_110001_10010; 
		2748: oled_colour = 16'b11111_110100_10010; 
		2749: oled_colour = 16'b11011_101011_10000; 
		2750: oled_colour = 16'b11010_100101_01110; 
		2825: oled_colour = 16'b01001_010100_00010; 
		2826: oled_colour = 16'b00101_010110_00010; 
		2827: oled_colour = 16'b00110_011000_00011; 
		2828: oled_colour = 16'b00110_010111_00011; 
		2829: oled_colour = 16'b01000_011011_00101; 
		2835: oled_colour = 16'b11101_110000_10010; 
		2836: oled_colour = 16'b11111_110101_10100; 
		2837: oled_colour = 16'b11110_101110_10001; 
		2838: oled_colour = 16'b11111_110110_10110; 
		2839: oled_colour = 16'b11111_110110_10111; 
		2840: oled_colour = 16'b11110_110000_10010; 
		2841: oled_colour = 16'b11100_101011_10000; 
		2842: oled_colour = 16'b11001_100100_01110; 
		2920: oled_colour = 16'b00101_011000_00100; 
		2921: oled_colour = 16'b10001_011110_01001; 
		2922: oled_colour = 16'b10010_010111_00110; 
		2923: oled_colour = 16'b10000_011010_00111; 
		2924: oled_colour = 16'b01110_010011_00011; 
		2925: oled_colour = 16'b10100_100001_01101; 
		2926: oled_colour = 16'b10011_100110_01111; 
		2934: oled_colour = 16'b11011_101010_01111; 
		3016: oled_colour = 16'b01101_011001_00111; 
		3017: oled_colour = 16'b10101_101000_01110; 
		3018: oled_colour = 16'b10001_011111_01010; 
		3019: oled_colour = 16'b11001_101100_10001; 
		3020: oled_colour = 16'b10111_100100_01101; 
		3021: oled_colour = 16'b01110_010111_00110; 
		3022: oled_colour = 16'b01001_011011_00111; 
		3023: oled_colour = 16'b10101_100000_01011; 
		3112: oled_colour = 16'b01101_100000_01001; 
		3113: oled_colour = 16'b10101_101111_10100; 
		3114: oled_colour = 16'b01101_101001_01110; 
		3115: oled_colour = 16'b11101_111110_11011; 
		3116: oled_colour = 16'b11011_110101_10110; 
		3117: oled_colour = 16'b01111_011111_01001; 
		3118: oled_colour = 16'b00111_010111_00100; 
		3119: oled_colour = 16'b10010_011100_01010; 
		3120: oled_colour = 16'b10110_110001_10010; 
		3121: oled_colour = 16'b11011_110011_10101; 
		3122: oled_colour = 16'b11100_101101_10011; 
		3208: oled_colour = 16'b10000_101100_01111; 
		3209: oled_colour = 16'b11000_110110_10111; 
		3210: oled_colour = 16'b11001_110110_10110; 
		3211: oled_colour = 16'b11100_110110_10110; 
		3212: oled_colour = 16'b11111_111100_11011; 
		3213: oled_colour = 16'b10111_110010_10100; 
		3214: oled_colour = 16'b01000_010111_00101; 
		3215: oled_colour = 16'b01110_011100_01001; 
		3216: oled_colour = 16'b11000_110110_10101; 
		3217: oled_colour = 16'b11111_111011_11001; 
		3218: oled_colour = 16'b11110_110100_10011; 
		3219: oled_colour = 16'b11111_101100_10001; 
		3220: oled_colour = 16'b11101_101001_10000; 
		3221: oled_colour = 16'b10101_100010_01100; 
		3305: oled_colour = 16'b11110_111001_11001; 
		3306: oled_colour = 16'b11111_110101_10111; 
		3307: oled_colour = 16'b11110_110000_10100; 
		3308: oled_colour = 16'b11111_110101_10110; 
		3309: oled_colour = 16'b11100_111011_10111; 
		3310: oled_colour = 16'b01100_100011_01010; 
		3311: oled_colour = 16'b01000_011010_00110; 
		3312: oled_colour = 16'b10000_101100_10001; 
		3313: oled_colour = 16'b10110_111000_10100; 
		3314: oled_colour = 16'b11010_110100_10011; 
		3315: oled_colour = 16'b11101_110011_10011; 
		3316: oled_colour = 16'b11000_110100_10010; 
		3317: oled_colour = 16'b11010_111011_10101; 
		3318: oled_colour = 16'b10100_110101_10010; 
		3401: oled_colour = 16'b11101_101111_10100; 
		3402: oled_colour = 16'b11110_111110_11011; 
		3403: oled_colour = 16'b10111_110000_10100; 
		3404: oled_colour = 16'b11011_110000_10000; 
		3405: oled_colour = 16'b11110_111000_10110; 
		3406: oled_colour = 16'b10000_101001_01110; 
		3408: oled_colour = 16'b10011_100100_01110; 
		3409: oled_colour = 16'b01110_100100_01101; 
		3410: oled_colour = 16'b01010_100000_01010; 
		3411: oled_colour = 16'b01101_100011_01011; 
		3412: oled_colour = 16'b01101_100111_01101; 
		3413: oled_colour = 16'b11001_111010_10100; 
		3414: oled_colour = 16'b11011_110111_10011; 
		3415: oled_colour = 16'b01011_011011_00111; 
		3498: oled_colour = 16'b10000_101100_01111; 
		3499: oled_colour = 16'b10011_110101_10100; 
		3500: oled_colour = 16'b11010_111011_10111; 
		3501: oled_colour = 16'b11111_111100_11100; 
		3502: oled_colour = 16'b10101_110000_10010; 
		3506: oled_colour = 16'b10000_011010_00111; 
		3507: oled_colour = 16'b11001_100101_01111; 
		3508: oled_colour = 16'b11001_111000_10100; 
		3509: oled_colour = 16'b11011_111110_10101; 
		3510: oled_colour = 16'b10011_101100_01111; 
		3593: oled_colour = 16'b10001_011000_00110; 
		3594: oled_colour = 16'b01001_010100_00011; 
		3595: oled_colour = 16'b10000_101011_01111; 
		3596: oled_colour = 16'b11110_111100_11101; 
		3598: oled_colour = 16'b10111_111001_10110; 
		3602: oled_colour = 16'b01100_100100_01100; 
		3603: oled_colour = 16'b11010_110111_10110; 
		3604: oled_colour = 16'b11111_111000_11001; 
		3605: oled_colour = 16'b11101_111000_10111; 
		3606: oled_colour = 16'b10001_100010_01100; 
		3688: oled_colour = 16'b10100_101000_01110; 
		3689: oled_colour = 16'b11111_111001_11010; 
		3690: oled_colour = 16'b11011_110100_10100; 
		3691: oled_colour = 16'b10100_101101_10000; 
		3692: oled_colour = 16'b11010_110110_10101; 
		3693: oled_colour = 16'b11101_111111_11011; 
		3694: oled_colour = 16'b10000_101100_10000; 
		3697: oled_colour = 16'b10010_011010_01000; 
		3698: oled_colour = 16'b01110_011101_01000; 
		3699: oled_colour = 16'b01010_100001_01010; 
		3700: oled_colour = 16'b01111_100011_01100; 
		3783: oled_colour = 16'b10100_100000_01010; 
		3784: oled_colour = 16'b01010_011010_00101; 
		3785: oled_colour = 16'b11100_110100_10101; 
		3786: oled_colour = 16'b11111_111100_11011; 
		3787: oled_colour = 16'b11110_110110_10101; 
		3788: oled_colour = 16'b10101_101111_10000; 
		3789: oled_colour = 16'b01110_101001_01110; 
		3793: oled_colour = 16'b01101_010010_00010; 
		3794: oled_colour = 16'b10011_011010_00111; 
		3795: oled_colour = 16'b10101_011111_01010; 
		3877: oled_colour = 16'b10000_010110_00100; 
		3878: oled_colour = 16'b01101_010010_00010; 
		3879: oled_colour = 16'b10111_100001_01100; 
		3880: oled_colour = 16'b01101_010111_00101; 
		3881: oled_colour = 16'b01100_011100_00111; 
		3889: oled_colour = 16'b01100_010001_00001; 
		3890: oled_colour = 16'b10011_011011_00111; 
		3972: oled_colour = 16'b10101_011100_01001; 
		3973: oled_colour = 16'b01100_010000_00001; 
		3974: oled_colour = 16'b10011_011011_00111; 
		3983: oled_colour = 16'b10111_100000_01100; 
		3984: oled_colour = 16'b10111_100000_01010; 
		3985: oled_colour = 16'b01011_010000_00001; 
		3986: oled_colour = 16'b10110_100000_01001; 
		4069: oled_colour = 16'b01100_010001_00001; 
		4070: oled_colour = 16'b10101_100001_01010; 
		4071: oled_colour = 16'b11001_100110_01110; 
		4080: oled_colour = 16'b10001_011000_00111; 
		4081: oled_colour = 16'b01100_010001_00010; 
		4082: oled_colour = 16'b10011_011001_00111; 
		4083: oled_colour = 16'b11001_100100_01110; 
		4165: oled_colour = 16'b10010_011000_00110; 
		4166: oled_colour = 16'b11011_101110_10010; 
		4167: oled_colour = 16'b11110_110010_10100; 
		4168: oled_colour = 16'b10101_011011_01010; 
		4179: oled_colour = 16'b11001_100011_01101; 
		4180: oled_colour = 16'b11011_101001_10001; 
		default: oled_colour = 16'b00000_000000_00000; 
	endcase
end

endmodule