module Gui_State2(
    input [12:0] pixel_index, 
    output reg [15:0] oled_colour 
); 

always@(pixel_index) 
begin
	case(pixel_index)
		1871: oled_colour = 16'b11111_111110_11111; 
		1872: oled_colour = 16'b11111_111001_11011; 
		1873: oled_colour = 16'b11111_111010_11100; 
		1874: oled_colour = 16'b11111_111110_11101; 
		1875: oled_colour = 16'b11111_111110_11010; 
		1876: oled_colour = 16'b11111_111110_11011; 
		1877: oled_colour = 16'b11111_111101_11011; 
		1878: oled_colour = 16'b11111_111101_11101; 
		1879: oled_colour = 16'b11111_111111_11110; 
		1880: oled_colour = 16'b11111_111111_11110; 
		1968: oled_colour = 16'b11111_111101_11101; 
		1969: oled_colour = 16'b11100_101101_01111; 
		1970: oled_colour = 16'b11101_110000_01100; 
		1971: oled_colour = 16'b11110_110110_01000; 
		1972: oled_colour = 16'b11101_110010_00111; 
		1973: oled_colour = 16'b11110_110100_01010; 
		1974: oled_colour = 16'b11101_110001_01000; 
		1975: oled_colour = 16'b11110_110110_10001; 
		1976: oled_colour = 16'b11111_111010_11010; 
		1977: oled_colour = 16'b11111_111110_11111; 
		2060: oled_colour = 16'b11111_111101_11110; 
		2061: oled_colour = 16'b11110_110101_11010; 
		2062: oled_colour = 16'b11101_110110_11001; 
		2063: oled_colour = 16'b10110_110001_10110; 
		2064: oled_colour = 16'b11001_110010_10111; 
		2065: oled_colour = 16'b11000_100110_10000; 
		2066: oled_colour = 16'b11100_101101_01011; 
		2067: oled_colour = 16'b11100_101110_01110; 
		2068: oled_colour = 16'b11101_110001_10010; 
		2069: oled_colour = 16'b11100_101110_01101; 
		2070: oled_colour = 16'b11110_110110_11000; 
		2155: oled_colour = 16'b11110_111100_11110; 
		2156: oled_colour = 16'b11001_101000_10001; 
		2157: oled_colour = 16'b11101_101111_10011; 
		2158: oled_colour = 16'b11111_111000_11001; 
		2159: oled_colour = 16'b10010_100001_01001; 
		2160: oled_colour = 16'b01000_010010_00001; 
		2161: oled_colour = 16'b10100_011100_01010; 
		2162: oled_colour = 16'b11001_100111_10000; 
		2163: oled_colour = 16'b11100_101011_10000; 
		2164: oled_colour = 16'b11010_101101_10101; 
		2165: oled_colour = 16'b11001_101000_10010; 
		2166: oled_colour = 16'b11100_110010_11000; 
		2168: oled_colour = 16'b11110_111000_11011; 
		2169: oled_colour = 16'b11111_111010_11101; 
		2251: oled_colour = 16'b10111_101110_10101; 
		2252: oled_colour = 16'b11001_100010_01100; 
		2253: oled_colour = 16'b11001_100110_10010; 
		2254: oled_colour = 16'b10101_101010_10111; 
		2255: oled_colour = 16'b11011_101000_01111; 
		2256: oled_colour = 16'b01100_011000_00110; 
		2257: oled_colour = 16'b11000_100011_01101; 
		2258: oled_colour = 16'b11000_100101_01110; 
		2259: oled_colour = 16'b11001_100111_01111; 
		2260: oled_colour = 16'b11100_101110_10100; 
		2261: oled_colour = 16'b11000_101001_01111; 
		2262: oled_colour = 16'b11010_101001_10000; 
		2263: oled_colour = 16'b11010_101101_10100; 
		2264: oled_colour = 16'b10110_011111_01011; 
		2265: oled_colour = 16'b10111_100010_01100; 
		2266: oled_colour = 16'b11101_110100_11001; 
		2347: oled_colour = 16'b10101_101110_10100; 
		2348: oled_colour = 16'b11000_100001_01011; 
		2349: oled_colour = 16'b11101_100011_01101; 
		2350: oled_colour = 16'b11100_110001_10110; 
		2351: oled_colour = 16'b11110_110110_11001; 
		2352: oled_colour = 16'b10100_011100_01001; 
		2353: oled_colour = 16'b11100_101100_10001; 
		2354: oled_colour = 16'b11110_101010_10001; 
		2355: oled_colour = 16'b11000_100011_01111; 
		2356: oled_colour = 16'b10100_100000_01011; 
		2357: oled_colour = 16'b10011_100000_01011; 
		2358: oled_colour = 16'b11010_100111_01111; 
		2359: oled_colour = 16'b11010_101011_10011; 
		2360: oled_colour = 16'b11000_100100_01110; 
		2361: oled_colour = 16'b11000_100011_01101; 
		2362: oled_colour = 16'b11001_101000_10001; 
		2443: oled_colour = 16'b10100_101110_10100; 
		2444: oled_colour = 16'b10000_011110_01000; 
		2445: oled_colour = 16'b11010_100101_01111; 
		2446: oled_colour = 16'b11010_100111_01110; 
		2447: oled_colour = 16'b11001_100101_01110; 
		2448: oled_colour = 16'b11100_101110_10011; 
		2449: oled_colour = 16'b11111_110110_10111; 
		2450: oled_colour = 16'b10100_011111_01010; 
		2451: oled_colour = 16'b01111_011010_01000; 
		2452: oled_colour = 16'b01010_011011_00111; 
		2453: oled_colour = 16'b01010_011100_01000; 
		2454: oled_colour = 16'b11010_101011_10010; 
		2455: oled_colour = 16'b10111_011111_01100; 
		2456: oled_colour = 16'b11011_101011_10010; 
		2457: oled_colour = 16'b11011_101101_10100; 
		2458: oled_colour = 16'b11110_111011_11101; 
		2539: oled_colour = 16'b11011_111001_11011; 
		2540: oled_colour = 16'b00100_010100_00001; 
		2541: oled_colour = 16'b10011_011001_01001; 
		2542: oled_colour = 16'b11000_100010_01110; 
		2543: oled_colour = 16'b11110_110111_11001; 
		2544: oled_colour = 16'b11111_111101_11110; 
		2545: oled_colour = 16'b10001_100000_01010; 
		2546: oled_colour = 16'b00101_011000_00100; 
		2547: oled_colour = 16'b01000_011101_01001; 
		2548: oled_colour = 16'b01001_011011_00111; 
		2549: oled_colour = 16'b10000_011010_01000; 
		2550: oled_colour = 16'b10111_011110_01011; 
		2551: oled_colour = 16'b11110_110011_10110; 
		2552: oled_colour = 16'b11011_101100_10011; 
		2553: oled_colour = 16'b11111_111100_11110; 
		2636: oled_colour = 16'b01011_100001_01010; 
		2637: oled_colour = 16'b01110_010111_00101; 
		2638: oled_colour = 16'b11110_101100_10011; 
		2639: oled_colour = 16'b11111_111000_11010; 
		2640: oled_colour = 16'b10110_100111_01111; 
		2641: oled_colour = 16'b00011_010011_00001; 
		2642: oled_colour = 16'b00111_011010_00101; 
		2643: oled_colour = 16'b10111_110011_10111; 
		2644: oled_colour = 16'b11011_110011_11000; 
		2645: oled_colour = 16'b10101_011001_01001; 
		2646: oled_colour = 16'b11100_101011_10001; 
		2647: oled_colour = 16'b11100_101101_10011; 
		2648: oled_colour = 16'b11100_110001_10111; 
		2732: oled_colour = 16'b10000_100110_01111; 
		2733: oled_colour = 16'b10000_011101_01001; 
		2734: oled_colour = 16'b10011_100001_01100; 
		2735: oled_colour = 16'b10011_011110_01011; 
		2736: oled_colour = 16'b10000_011000_00110; 
		2737: oled_colour = 16'b01110_011111_01010; 
		2738: oled_colour = 16'b10001_011110_01010; 
		2741: oled_colour = 16'b11011_110001_10111; 
		2742: oled_colour = 16'b11011_101010_10010; 
		2743: oled_colour = 16'b11011_110000_10111; 
		2827: oled_colour = 16'b11101_111001_11100; 
		2828: oled_colour = 16'b01110_010101_00101; 
		2829: oled_colour = 16'b10110_100010_01101; 
		2830: oled_colour = 16'b10101_100110_01110; 
		2831: oled_colour = 16'b10011_100101_01100; 
		2832: oled_colour = 16'b01110_010101_00101; 
		2833: oled_colour = 16'b01000_011100_00110; 
		2834: oled_colour = 16'b10010_011101_01001; 
		2835: oled_colour = 16'b11101_111000_11100; 
		2923: oled_colour = 16'b11011_111001_11010; 
		2924: oled_colour = 16'b10000_100110_01101; 
		2925: oled_colour = 16'b10000_100111_01111; 
		2926: oled_colour = 16'b11100_111000_10100; 
		2927: oled_colour = 16'b10101_101010_01111; 
		2928: oled_colour = 16'b01100_011010_00111; 
		2929: oled_colour = 16'b01010_011101_00111; 
		2930: oled_colour = 16'b01110_011101_01001; 
		2931: oled_colour = 16'b10101_101111_10110; 
		3019: oled_colour = 16'b11011_111001_11011; 
		3020: oled_colour = 16'b10010_101110_10010; 
		3021: oled_colour = 16'b10011_101111_10100; 
		3022: oled_colour = 16'b11001_110011_10010; 
		3023: oled_colour = 16'b11011_110000_10010; 
		3024: oled_colour = 16'b10010_101000_01110; 
		3025: oled_colour = 16'b00111_011011_00101; 
		3026: oled_colour = 16'b01110_011110_01010; 
		3027: oled_colour = 16'b10001_100001_01100; 
		3028: oled_colour = 16'b11010_110011_11000; 
		3115: oled_colour = 16'b11111_111110_11110; 
		3116: oled_colour = 16'b11000_110000_10010; 
		3117: oled_colour = 16'b11011_110101_11000; 
		3118: oled_colour = 16'b11100_110001_10110; 
		3119: oled_colour = 16'b11110_110010_10110; 
		3120: oled_colour = 16'b10111_101001_10001; 
		3121: oled_colour = 16'b00111_010110_00100; 
		3122: oled_colour = 16'b10011_100000_01100; 
		3123: oled_colour = 16'b11111_110010_10110; 
		3124: oled_colour = 16'b11011_101101_10010; 
		3125: oled_colour = 16'b11101_110111_11011; 
		3212: oled_colour = 16'b11101_110011_10101; 
		3213: oled_colour = 16'b11101_111010_11001; 
		3214: oled_colour = 16'b11011_101111_10100; 
		3215: oled_colour = 16'b11111_101101_10001; 
		3216: oled_colour = 16'b10111_110001_10011; 
		3217: oled_colour = 16'b01000_011110_01001; 
		3218: oled_colour = 16'b01100_100000_01011; 
		3219: oled_colour = 16'b10101_110011_10100; 
		3220: oled_colour = 16'b11101_111000_10110; 
		3221: oled_colour = 16'b10111_100000_01011; 
		3222: oled_colour = 16'b11010_101111_10111; 
		3308: oled_colour = 16'b11010_111000_11001; 
		3309: oled_colour = 16'b10000_101011_01111; 
		3310: oled_colour = 16'b10011_101100_10001; 
		3311: oled_colour = 16'b11100_110101_10010; 
		3312: oled_colour = 16'b11101_110000_10010; 
		3313: oled_colour = 16'b01101_011100_01000; 
		3314: oled_colour = 16'b01001_011110_01001; 
		3315: oled_colour = 16'b10001_101100_10010; 
		3316: oled_colour = 16'b11001_110011_10011; 
		3317: oled_colour = 16'b11111_110111_10111; 
		3318: oled_colour = 16'b10100_100111_01111; 
		3319: oled_colour = 16'b11010_110110_11010; 
		3405: oled_colour = 16'b01101_100011_01101; 
		3406: oled_colour = 16'b01000_011101_01000; 
		3407: oled_colour = 16'b10101_110111_10100; 
		3408: oled_colour = 16'b11100_111110_10101; 
		3409: oled_colour = 16'b01111_100011_01100; 
		3410: oled_colour = 16'b10001_100010_01011; 
		3411: oled_colour = 16'b01101_100100_01101; 
		3412: oled_colour = 16'b01110_101000_01110; 
		3413: oled_colour = 16'b11000_111010_11000; 
		3414: oled_colour = 16'b10101_101110_10001; 
		3415: oled_colour = 16'b01111_100000_01011; 
		3501: oled_colour = 16'b10100_100110_01111; 
		3502: oled_colour = 16'b01001_010011_00011; 
		3503: oled_colour = 16'b10100_101011_10000; 
		3504: oled_colour = 16'b10111_111010_10100; 
		3505: oled_colour = 16'b01111_101010_10000; 
		3506: oled_colour = 16'b11010_110101_11001; 
		3507: oled_colour = 16'b01001_011001_00110; 
		3508: oled_colour = 16'b01001_011101_01001; 
		3509: oled_colour = 16'b10000_110000_10010; 
		3510: oled_colour = 16'b10010_101111_10001; 
		3511: oled_colour = 16'b10000_100001_01100; 
		3512: oled_colour = 16'b11111_111100_11110; 
		3596: oled_colour = 16'b11010_110100_11000; 
		3597: oled_colour = 16'b11000_101001_01111; 
		3598: oled_colour = 16'b10000_100011_01101; 
		3599: oled_colour = 16'b01111_101000_10000; 
		3600: oled_colour = 16'b01110_100010_01100; 
		3601: oled_colour = 16'b10010_101000_10001; 
		3603: oled_colour = 16'b10111_101010_10011; 
		3604: oled_colour = 16'b01110_011000_00111; 
		3605: oled_colour = 16'b11001_101100_10011; 
		3606: oled_colour = 16'b11011_110111_10111; 
		3607: oled_colour = 16'b11000_101011_10001; 
		3608: oled_colour = 16'b11111_111100_11110; 
		3692: oled_colour = 16'b10111_101011_10011; 
		3693: oled_colour = 16'b01100_011011_00111; 
		3694: oled_colour = 16'b11000_101100_10010; 
		3695: oled_colour = 16'b10111_101001_10010; 
		3696: oled_colour = 16'b01111_011011_01001; 
		3697: oled_colour = 16'b11101_111001_11100; 
		3699: oled_colour = 16'b11110_111101_11110; 
		3700: oled_colour = 16'b01101_100000_01011; 
		3701: oled_colour = 16'b01111_011011_01000; 
		3702: oled_colour = 16'b01111_100101_01101; 
		3703: oled_colour = 16'b01101_011110_01001; 
		3704: oled_colour = 16'b11110_111100_11110; 
		3788: oled_colour = 16'b11101_110101_11001; 
		3789: oled_colour = 16'b10010_011010_00111; 
		3790: oled_colour = 16'b01101_011010_00111; 
		3791: oled_colour = 16'b01011_011001_00110; 
		3792: oled_colour = 16'b11000_110100_11000; 
		3796: oled_colour = 16'b11101_111100_11101; 
		3797: oled_colour = 16'b01111_011101_01001; 
		3798: oled_colour = 16'b10010_011100_01000; 
		3799: oled_colour = 16'b10101_011111_01011; 
		3884: oled_colour = 16'b11101_110111_11011; 
		3885: oled_colour = 16'b10010_011001_00111; 
		3886: oled_colour = 16'b10010_011000_00110; 
		3887: oled_colour = 16'b10111_101000_10001; 
		3893: oled_colour = 16'b11011_110011_11000; 
		3894: oled_colour = 16'b01011_001110_00001; 
		3895: oled_colour = 16'b10001_011000_00110; 
		3896: oled_colour = 16'b11101_110101_11001; 
		3980: oled_colour = 16'b11010_101100_10100; 
		3981: oled_colour = 16'b01110_010010_00011; 
		3982: oled_colour = 16'b10000_010110_00101; 
		3983: oled_colour = 16'b11011_110011_11000; 
		3989: oled_colour = 16'b11100_110000_10110; 
		3990: oled_colour = 16'b10101_011110_01001; 
		3991: oled_colour = 16'b01100_010001_00001; 
		3992: oled_colour = 16'b10010_011001_00110; 
		3993: oled_colour = 16'b11100_110011_11000; 
		4076: oled_colour = 16'b11101_110100_11001; 
		4077: oled_colour = 16'b01111_010011_00011; 
		4078: oled_colour = 16'b10001_010101_00110; 
		4079: oled_colour = 16'b11011_101110_10100; 
		4080: oled_colour = 16'b11111_111101_11111; 
		4085: oled_colour = 16'b11101_110101_11000; 
		4086: oled_colour = 16'b11100_101100_10011; 
		4087: oled_colour = 16'b01111_010100_00011; 
		4088: oled_colour = 16'b01011_001110_00001; 
		4089: oled_colour = 16'b10101_011100_01001; 
		4090: oled_colour = 16'b11100_110000_10101; 
		4091: oled_colour = 16'b11101_110111_11011; 
		4173: oled_colour = 16'b11001_101011_10100; 
		4174: oled_colour = 16'b10111_100010_01101; 
		4175: oled_colour = 16'b11011_101010_10001; 
		4176: oled_colour = 16'b11010_101101_10101; 
		4183: oled_colour = 16'b11101_110101_11001; 
		4184: oled_colour = 16'b10111_100110_10000; 
		4185: oled_colour = 16'b11010_101010_10010; 
		4186: oled_colour = 16'b11010_101100_10011; 
		4187: oled_colour = 16'b11100_110000_10111; 
		default: oled_colour = 16'b00000_000000_00000; 
	endcase
end

endmodule