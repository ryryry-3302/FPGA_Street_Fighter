module Gui_State3(
    input [12:0] pixel_index, 
    output reg [15:0] oled_colour 
); 

always@(pixel_index) 
begin
	case(pixel_index)
		1680: oled_colour = 16'b11111_111111_11111; 
		1681: oled_colour = 16'b11111_111111_11111; 
		1682: oled_colour = 16'b11111_111111_11111; 
		1683: oled_colour = 16'b11111_111111_11111; 
		1684: oled_colour = 16'b11111_111111_11111; 
		1685: oled_colour = 16'b11111_111111_11111; 
		1686: oled_colour = 16'b11111_111111_11111; 
		1687: oled_colour = 16'b11111_111111_11111; 
		1688: oled_colour = 16'b11111_111111_11111; 
		1689: oled_colour = 16'b11111_111111_11111; 
		1868: oled_colour = 16'b11111_111111_11111; 
		1869: oled_colour = 16'b11111_111111_11111; 
		1870: oled_colour = 16'b11111_111111_11111; 
		1871: oled_colour = 16'b11111_111111_11111; 
		1872: oled_colour = 16'b11111_111010_11100; 
		1873: oled_colour = 16'b11110_110100_10111; 
		1874: oled_colour = 16'b11111_111000_11000; 
		1875: oled_colour = 16'b11111_111011_10110; 
		1876: oled_colour = 16'b11111_111100_10011; 
		1877: oled_colour = 16'b11111_111010_10110; 
		1878: oled_colour = 16'b11111_111011_10110; 
		1879: oled_colour = 16'b11111_111011_11000; 
		1880: oled_colour = 16'b11111_111100_11011; 
		1881: oled_colour = 16'b11111_111101_11110; 
		1969: oled_colour = 16'b11110_111000_11001; 
		1970: oled_colour = 16'b11011_101010_01010; 
		1971: oled_colour = 16'b11110_110011_01010; 
		1972: oled_colour = 16'b11101_110010_00110; 
		1973: oled_colour = 16'b11110_110010_01001; 
		1974: oled_colour = 16'b11110_110010_01000; 
		1975: oled_colour = 16'b11110_110100_01110; 
		1976: oled_colour = 16'b11111_111011_11001; 
		1977: oled_colour = 16'b11111_111110_11110; 
		1978: oled_colour = 16'b11111_111111_11111; 
		2058: oled_colour = 16'b11111_111111_11111; 
		2060: oled_colour = 16'b11111_111110_11111; 
		2061: oled_colour = 16'b11100_101111_10110; 
		2062: oled_colour = 16'b11111_110100_10111; 
		2063: oled_colour = 16'b10111_101110_10011; 
		2064: oled_colour = 16'b10001_100111_01111; 
		2065: oled_colour = 16'b10101_100100_01111; 
		2066: oled_colour = 16'b11000_100101_01110; 
		2067: oled_colour = 16'b11101_101111_01100; 
		2068: oled_colour = 16'b11011_101101_10011; 
		2069: oled_colour = 16'b11100_110001_10010; 
		2070: oled_colour = 16'b11101_101111_10011; 
		2075: oled_colour = 16'b11111_111111_11111; 
		2154: oled_colour = 16'b11111_111111_11111; 
		2155: oled_colour = 16'b11111_111111_11111; 
		2156: oled_colour = 16'b11000_101010_10011; 
		2157: oled_colour = 16'b11011_101010_10000; 
		2158: oled_colour = 16'b11100_110110_11001; 
		2159: oled_colour = 16'b11101_110001_10101; 
		2160: oled_colour = 16'b01010_010101_00010; 
		2161: oled_colour = 16'b01110_010111_00101; 
		2162: oled_colour = 16'b10110_100010_01110; 
		2163: oled_colour = 16'b11010_101000_01111; 
		2164: oled_colour = 16'b11100_101110_10011; 
		2165: oled_colour = 16'b11001_101001_10011; 
		2166: oled_colour = 16'b11010_101011_10010; 
		2167: oled_colour = 16'b11110_111000_11011; 
		2168: oled_colour = 16'b11101_110110_11010; 
		2169: oled_colour = 16'b11011_101111_10101; 
		2170: oled_colour = 16'b11111_111011_11101; 
		2172: oled_colour = 16'b11111_111111_11111; 
		2249: oled_colour = 16'b11111_111111_11111; 
		2251: oled_colour = 16'b11110_111110_11111; 
		2252: oled_colour = 16'b10011_100000_01011; 
		2253: oled_colour = 16'b11110_100101_01110; 
		2254: oled_colour = 16'b10011_011111_10001; 
		2255: oled_colour = 16'b11100_110000_10111; 
		2256: oled_colour = 16'b10100_011111_01011; 
		2257: oled_colour = 16'b10010_011111_01010; 
		2258: oled_colour = 16'b11100_101000_01111; 
		2259: oled_colour = 16'b11000_100101_01110; 
		2260: oled_colour = 16'b11011_101010_10001; 
		2261: oled_colour = 16'b11001_101001_10000; 
		2262: oled_colour = 16'b11001_100111_01110; 
		2263: oled_colour = 16'b11001_101000_10001; 
		2264: oled_colour = 16'b11001_101000_10000; 
		2265: oled_colour = 16'b10101_011011_01001; 
		2266: oled_colour = 16'b11001_100110_01110; 
		2267: oled_colour = 16'b11111_111010_11100; 
		2269: oled_colour = 16'b11111_111111_11111; 
		2345: oled_colour = 16'b11111_111111_11111; 
		2347: oled_colour = 16'b11110_111110_11111; 
		2348: oled_colour = 16'b10000_100000_01010; 
		2349: oled_colour = 16'b11110_100111_01111; 
		2350: oled_colour = 16'b11101_101010_01111; 
		2351: oled_colour = 16'b11111_111011_11011; 
		2352: oled_colour = 16'b11000_100011_01110; 
		2353: oled_colour = 16'b11001_100111_01110; 
		2354: oled_colour = 16'b11111_101101_10010; 
		2355: oled_colour = 16'b11010_100100_01111; 
		2356: oled_colour = 16'b10100_011110_01011; 
		2357: oled_colour = 16'b01111_011100_01000; 
		2358: oled_colour = 16'b10110_100100_01101; 
		2359: oled_colour = 16'b11011_101100_10011; 
		2360: oled_colour = 16'b11000_100100_01111; 
		2361: oled_colour = 16'b11010_100111_10000; 
		2362: oled_colour = 16'b11000_100100_01110; 
		2363: oled_colour = 16'b11110_111000_11100; 
		2365: oled_colour = 16'b11111_111111_11111; 
		2441: oled_colour = 16'b11111_111111_11111; 
		2442: oled_colour = 16'b11111_111111_11111; 
		2443: oled_colour = 16'b11111_111111_11111; 
		2444: oled_colour = 16'b01011_011110_01000; 
		2445: oled_colour = 16'b10101_011111_01011; 
		2446: oled_colour = 16'b10111_100000_01100; 
		2447: oled_colour = 16'b11001_100101_01101; 
		2448: oled_colour = 16'b11011_101100_10010; 
		2449: oled_colour = 16'b11111_111010_11010; 
		2450: oled_colour = 16'b10110_100101_01101; 
		2451: oled_colour = 16'b01101_011001_00111; 
		2452: oled_colour = 16'b01011_011011_00111; 
		2453: oled_colour = 16'b00111_011010_00110; 
		2454: oled_colour = 16'b10011_100011_01100; 
		2455: oled_colour = 16'b11000_100010_01110; 
		2456: oled_colour = 16'b11010_101000_10000; 
		2457: oled_colour = 16'b11100_101110_10100; 
		2458: oled_colour = 16'b11110_111001_11100; 
		2460: oled_colour = 16'b11111_111111_11111; 
		2538: oled_colour = 16'b11111_111111_11111; 
		2540: oled_colour = 16'b01110_100111_01110; 
		2541: oled_colour = 16'b01000_010011_00010; 
		2542: oled_colour = 16'b11000_011101_01100; 
		2543: oled_colour = 16'b11101_110010_10110; 
		2544: oled_colour = 16'b11111_111111_11111; 
		2545: oled_colour = 16'b10111_101001_10001; 
		2546: oled_colour = 16'b00100_010011_00001; 
		2547: oled_colour = 16'b00111_011100_01000; 
		2548: oled_colour = 16'b01011_100001_01011; 
		2549: oled_colour = 16'b01111_011010_01000; 
		2550: oled_colour = 16'b10101_011010_01001; 
		2551: oled_colour = 16'b11101_101111_10100; 
		2552: oled_colour = 16'b11100_110001_10101; 
		2553: oled_colour = 16'b11101_110101_11001; 
		2555: oled_colour = 16'b11111_111111_11111; 
		2634: oled_colour = 16'b11111_111111_11111; 
		2636: oled_colour = 16'b11001_110101_11001; 
		2637: oled_colour = 16'b00111_010011_00010; 
		2638: oled_colour = 16'b11000_100110_01111; 
		2639: oled_colour = 16'b11110_110000_10100; 
		2640: oled_colour = 16'b10111_101000_10000; 
		2641: oled_colour = 16'b00101_010100_00001; 
		2642: oled_colour = 16'b00010_010100_00001; 
		2643: oled_colour = 16'b10101_101110_10100; 
		2644: oled_colour = 16'b11111_111110_11111; 
		2645: oled_colour = 16'b11001_101001_10011; 
		2646: oled_colour = 16'b11001_100000_01011; 
		2647: oled_colour = 16'b11101_101111_10011; 
		2648: oled_colour = 16'b11001_101010_10011; 
		2649: oled_colour = 16'b11111_111111_11111; 
		2650: oled_colour = 16'b11111_111111_11111; 
		2730: oled_colour = 16'b11111_111111_11111; 
		2732: oled_colour = 16'b10101_101100_10010; 
		2733: oled_colour = 16'b01010_011001_00110; 
		2734: oled_colour = 16'b10000_011001_00111; 
		2735: oled_colour = 16'b10100_011101_01010; 
		2736: oled_colour = 16'b01110_011010_00111; 
		2737: oled_colour = 16'b01111_100100_01101; 
		2738: oled_colour = 16'b01101_011000_00110; 
		2739: oled_colour = 16'b11001_110101_11000; 
		2741: oled_colour = 16'b11111_111111_11111; 
		2742: oled_colour = 16'b11110_110101_11001; 
		2743: oled_colour = 16'b11110_111000_11011; 
		2744: oled_colour = 16'b11111_111111_11111; 
		2825: oled_colour = 16'b11111_111111_11111; 
		2827: oled_colour = 16'b11101_111010_11100; 
		2828: oled_colour = 16'b10001_011111_01011; 
		2829: oled_colour = 16'b10101_100011_01101; 
		2830: oled_colour = 16'b10010_011001_01000; 
		2831: oled_colour = 16'b10001_011011_01000; 
		2832: oled_colour = 16'b10000_101010_01111; 
		2833: oled_colour = 16'b01010_011110_01000; 
		2834: oled_colour = 16'b10001_011010_00111; 
		2835: oled_colour = 16'b11010_110010_10111; 
		2836: oled_colour = 16'b11111_111111_11111; 
		2837: oled_colour = 16'b11111_111111_11111; 
		2921: oled_colour = 16'b11111_111111_11111; 
		2923: oled_colour = 16'b11101_111100_11101; 
		2924: oled_colour = 16'b10001_101011_10000; 
		2925: oled_colour = 16'b10011_101011_10001; 
		2926: oled_colour = 16'b10101_101000_01111; 
		2927: oled_colour = 16'b10000_011011_00111; 
		2928: oled_colour = 16'b01001_011101_00111; 
		2929: oled_colour = 16'b01001_011010_00101; 
		2930: oled_colour = 16'b10110_100111_01110; 
		2931: oled_colour = 16'b10101_101110_10011; 
		2933: oled_colour = 16'b11111_111111_11111; 
		2934: oled_colour = 16'b11111_111111_11111; 
		2935: oled_colour = 16'b11111_111111_11111; 
		3017: oled_colour = 16'b11111_111111_11111; 
		3018: oled_colour = 16'b11111_111111_11111; 
		3019: oled_colour = 16'b11011_111010_11011; 
		3020: oled_colour = 16'b10110_110010_10110; 
		3021: oled_colour = 16'b10101_110101_10100; 
		3022: oled_colour = 16'b10100_110110_10010; 
		3023: oled_colour = 16'b01101_100111_01101; 
		3024: oled_colour = 16'b00111_011001_00110; 
		3025: oled_colour = 16'b00111_010111_00100; 
		3026: oled_colour = 16'b01110_101001_01110; 
		3027: oled_colour = 16'b10001_101101_10010; 
		3028: oled_colour = 16'b11110_111101_11110; 
		3030: oled_colour = 16'b11111_111111_11111; 
		3114: oled_colour = 16'b11111_111111_11111; 
		3115: oled_colour = 16'b10110_110010_10101; 
		3116: oled_colour = 16'b11000_110010_10010; 
		3117: oled_colour = 16'b11100_101111_10010; 
		3118: oled_colour = 16'b11111_110111_10100; 
		3119: oled_colour = 16'b10111_110011_10011; 
		3120: oled_colour = 16'b01000_011000_00101; 
		3121: oled_colour = 16'b01110_011010_01000; 
		3122: oled_colour = 16'b10110_101110_10001; 
		3123: oled_colour = 16'b11010_101110_10010; 
		3124: oled_colour = 16'b11101_110100_11000; 
		3125: oled_colour = 16'b11111_111111_11111; 
		3126: oled_colour = 16'b11111_111111_11111; 
		3209: oled_colour = 16'b11111_111111_11111; 
		3210: oled_colour = 16'b11111_111111_11111; 
		3211: oled_colour = 16'b11100_110010_10101; 
		3212: oled_colour = 16'b11110_110100_10110; 
		3213: oled_colour = 16'b11110_110101_11000; 
		3214: oled_colour = 16'b11110_111010_11011; 
		3215: oled_colour = 16'b11001_110100_10101; 
		3216: oled_colour = 16'b01000_011001_00110; 
		3217: oled_colour = 16'b01110_100011_01100; 
		3218: oled_colour = 16'b11101_110111_10110; 
		3219: oled_colour = 16'b11110_111000_11000; 
		3220: oled_colour = 16'b11100_101111_10100; 
		3221: oled_colour = 16'b11111_111110_11111; 
		3223: oled_colour = 16'b11111_111111_11111; 
		3304: oled_colour = 16'b11111_111111_11111; 
		3307: oled_colour = 16'b11010_110100_10111; 
		3308: oled_colour = 16'b11100_110010_10111; 
		3309: oled_colour = 16'b11101_101110_10010; 
		3310: oled_colour = 16'b11111_111101_11011; 
		3311: oled_colour = 16'b10101_110011_10010; 
		3312: oled_colour = 16'b00101_010111_00100; 
		3313: oled_colour = 16'b10001_101011_10001; 
		3314: oled_colour = 16'b11001_110111_10100; 
		3315: oled_colour = 16'b11110_111000_10101; 
		3316: oled_colour = 16'b11100_101010_10000; 
		3317: oled_colour = 16'b11100_110001_11000; 
		3319: oled_colour = 16'b11111_111111_11111; 
		3399: oled_colour = 16'b11111_111111_11111; 
		3401: oled_colour = 16'b11111_111111_11111; 
		3402: oled_colour = 16'b11100_110010_10111; 
		3403: oled_colour = 16'b10100_100100_01101; 
		3404: oled_colour = 16'b10000_011111_01001; 
		3405: oled_colour = 16'b11000_100110_01110; 
		3406: oled_colour = 16'b11110_110011_10110; 
		3407: oled_colour = 16'b10100_101010_10000; 
		3408: oled_colour = 16'b01111_100000_01100; 
		3409: oled_colour = 16'b01110_100000_01010; 
		3410: oled_colour = 16'b01111_101110_10000; 
		3411: oled_colour = 16'b11010_110111_10110; 
		3412: oled_colour = 16'b10111_101111_10010; 
		3413: oled_colour = 16'b10101_100110_01110; 
		3414: oled_colour = 16'b11111_111111_11111; 
		3494: oled_colour = 16'b11111_111111_11111; 
		3495: oled_colour = 16'b11111_111111_11111; 
		3496: oled_colour = 16'b11100_111001_11100; 
		3497: oled_colour = 16'b10000_011100_01001; 
		3498: oled_colour = 16'b10110_101010_01111; 
		3499: oled_colour = 16'b10111_100100_01110; 
		3500: oled_colour = 16'b10010_110011_10001; 
		3501: oled_colour = 16'b11001_111010_10100; 
		3502: oled_colour = 16'b11000_110110_10101; 
		3503: oled_colour = 16'b01111_101011_10000; 
		3504: oled_colour = 16'b10011_100011_01111; 
		3505: oled_colour = 16'b10000_011000_00111; 
		3506: oled_colour = 16'b10111_110001_10011; 
		3507: oled_colour = 16'b10011_110101_10100; 
		3508: oled_colour = 16'b01101_100001_01010; 
		3509: oled_colour = 16'b10100_101000_10001; 
		3511: oled_colour = 16'b11111_111111_11111; 
		3589: oled_colour = 16'b11111_111111_11111; 
		3590: oled_colour = 16'b11111_111111_11111; 
		3592: oled_colour = 16'b10011_100011_01101; 
		3593: oled_colour = 16'b01100_011101_00111; 
		3594: oled_colour = 16'b11101_111011_11000; 
		3595: oled_colour = 16'b11111_110110_11000; 
		3596: oled_colour = 16'b11000_110001_10011; 
		3597: oled_colour = 16'b10100_101111_10001; 
		3598: oled_colour = 16'b01110_101001_01101; 
		3599: oled_colour = 16'b10111_110010_10111; 
		3600: oled_colour = 16'b10001_100101_01111; 
		3601: oled_colour = 16'b10000_100010_01100; 
		3602: oled_colour = 16'b11010_101011_10010; 
		3603: oled_colour = 16'b10111_101011_10001; 
		3604: oled_colour = 16'b11001_101100_10011; 
		3605: oled_colour = 16'b11111_111111_11111; 
		3606: oled_colour = 16'b11111_111111_11111; 
		3607: oled_colour = 16'b11111_111111_11111; 
		3685: oled_colour = 16'b11111_111111_11111; 
		3686: oled_colour = 16'b11111_111111_11111; 
		3687: oled_colour = 16'b10101_100101_01111; 
		3688: oled_colour = 16'b10101_011101_01001; 
		3689: oled_colour = 16'b10000_011100_01000; 
		3690: oled_colour = 16'b01100_100001_01001; 
		3691: oled_colour = 16'b10010_101010_01111; 
		3692: oled_colour = 16'b10111_101110_10100; 
		3693: oled_colour = 16'b11100_110001_10111; 
		3694: oled_colour = 16'b11100_111000_11011; 
		3695: oled_colour = 16'b11111_111110_11111; 
		3696: oled_colour = 16'b10101_100010_01100; 
		3697: oled_colour = 16'b01110_100010_01010; 
		3698: oled_colour = 16'b01001_011101_01000; 
		3699: oled_colour = 16'b10101_101100_10011; 
		3701: oled_colour = 16'b11111_111111_11111; 
		3778: oled_colour = 16'b11111_111111_11111; 
		3780: oled_colour = 16'b11111_111100_11110; 
		3781: oled_colour = 16'b11101_101111_10101; 
		3782: oled_colour = 16'b11001_101000_10001; 
		3783: oled_colour = 16'b01101_010001_00010; 
		3784: oled_colour = 16'b10000_010100_00100; 
		3785: oled_colour = 16'b10101_011110_01011; 
		3786: oled_colour = 16'b10110_101010_10010; 
		3787: oled_colour = 16'b11010_110111_11010; 
		3788: oled_colour = 16'b11110_111110_11111; 
		3791: oled_colour = 16'b10110_100111_10000; 
		3792: oled_colour = 16'b01111_010100_00100; 
		3793: oled_colour = 16'b10111_100000_01011; 
		3794: oled_colour = 16'b11001_101110_10101; 
		3796: oled_colour = 16'b11111_111111_11111; 
		3797: oled_colour = 16'b11111_111111_11111; 
		3874: oled_colour = 16'b11111_111111_11111; 
		3876: oled_colour = 16'b11111_111100_11110; 
		3877: oled_colour = 16'b10111_011111_01011; 
		3878: oled_colour = 16'b10000_010101_00100; 
		3879: oled_colour = 16'b10010_011010_01000; 
		3880: oled_colour = 16'b11011_110000_10110; 
		3881: oled_colour = 16'b11111_111111_11111; 
		3885: oled_colour = 16'b11111_111111_11111; 
		3886: oled_colour = 16'b11011_101110_10101; 
		3887: oled_colour = 16'b10010_011000_00111; 
		3888: oled_colour = 16'b01111_010110_00100; 
		3889: oled_colour = 16'b10111_100101_01111; 
		3891: oled_colour = 16'b11111_111111_11111; 
		3973: oled_colour = 16'b10000_011010_00111; 
		3974: oled_colour = 16'b01100_001111_00001; 
		3975: oled_colour = 16'b10110_100011_01110; 
		3978: oled_colour = 16'b11111_111111_11111; 
		3979: oled_colour = 16'b11111_111111_11111; 
		3980: oled_colour = 16'b11111_111111_11111; 
		3982: oled_colour = 16'b11011_101101_10100; 
		3983: oled_colour = 16'b01111_010011_00100; 
		3984: oled_colour = 16'b01101_010011_00010; 
		3985: oled_colour = 16'b10111_100100_01101; 
		3986: oled_colour = 16'b11111_111111_11111; 
		3988: oled_colour = 16'b11111_111111_11111; 
		4069: oled_colour = 16'b10101_011110_01011; 
		4070: oled_colour = 16'b11001_100011_01101; 
		4071: oled_colour = 16'b11001_100110_10000; 
		4072: oled_colour = 16'b11111_111100_11110; 
		4073: oled_colour = 16'b11111_111111_11111; 
		4074: oled_colour = 16'b11111_111111_11111; 
		4077: oled_colour = 16'b11111_111111_11111; 
		4079: oled_colour = 16'b11001_101101_10100; 
		4080: oled_colour = 16'b10001_010101_00101; 
		4081: oled_colour = 16'b10111_100000_01100; 
		4082: oled_colour = 16'b11011_101110_10101; 
		4083: oled_colour = 16'b11111_111100_11110; 
		4084: oled_colour = 16'b11111_111111_11111; 
		4085: oled_colour = 16'b11111_111111_11111; 
		4163: oled_colour = 16'b11111_111111_11111; 
		4165: oled_colour = 16'b11101_110101_11010; 
		4166: oled_colour = 16'b11000_100100_01111; 
		4167: oled_colour = 16'b11000_101000_10001; 
		4168: oled_colour = 16'b11111_111101_11110; 
		4170: oled_colour = 16'b11111_111111_11111; 
		4174: oled_colour = 16'b11111_111111_11111; 
		4176: oled_colour = 16'b11100_110010_11000; 
		4177: oled_colour = 16'b10111_100100_01111; 
		4178: oled_colour = 16'b10111_100100_01111; 
		4179: oled_colour = 16'b11101_110101_11010; 
		4181: oled_colour = 16'b11111_111111_11111; 
		4262: oled_colour = 16'b11111_111111_11111; 
		4263: oled_colour = 16'b11111_111111_11111; 
		4271: oled_colour = 16'b11111_111111_11111; 
		4273: oled_colour = 16'b11111_111111_11111; 
		4274: oled_colour = 16'b11111_111111_11111; 
		4357: oled_colour = 16'b11111_111111_11111; 
		4368: oled_colour = 16'b11111_111111_11111; 
		default: oled_colour = 16'b00000_000000_00000; 
	endcase
end

endmodule