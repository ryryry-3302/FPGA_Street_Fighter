module Gui_Inj1(
    input [12:0] pixel_index, 
    output reg [15:0] oled_colour 
); 

always@(pixel_index) 
begin
	case(pixel_index)
		2249: oled_colour = 16'b11111_111110_11111; 
		2250: oled_colour = 16'b11110_111000_11101; 
		2251: oled_colour = 16'b11011_110110_11011; 
		2252: oled_colour = 16'b10100_101101_10101; 
		2253: oled_colour = 16'b10100_101101_10101; 
		2254: oled_colour = 16'b11001_110110_11011; 
		2255: oled_colour = 16'b11110_111110_11111; 
		2342: oled_colour = 16'b11111_111110_11111; 
		2343: oled_colour = 16'b11110_111000_11101; 
		2344: oled_colour = 16'b11011_101110_10110; 
		2345: oled_colour = 16'b11010_100110_10000; 
		2346: oled_colour = 16'b11101_101110_10011; 
		2347: oled_colour = 16'b10111_100110_01110; 
		2348: oled_colour = 16'b00100_010100_00010; 
		2349: oled_colour = 16'b00010_010011_00001; 
		2350: oled_colour = 16'b01110_011101_01000; 
		2351: oled_colour = 16'b10110_100101_01110; 
		2352: oled_colour = 16'b01100_011111_01011; 
		2353: oled_colour = 16'b10110_101100_10100; 
		2354: oled_colour = 16'b11100_101111_10111; 
		2355: oled_colour = 16'b11110_110111_11010; 
		2356: oled_colour = 16'b11110_111000_11100; 
		2357: oled_colour = 16'b11111_111101_11111; 
		2437: oled_colour = 16'b11011_110010_11001; 
		2438: oled_colour = 16'b11011_101101_10101; 
		2439: oled_colour = 16'b11100_101100_10001; 
		2440: oled_colour = 16'b11011_011100_01000; 
		2441: oled_colour = 16'b11100_101101_10010; 
		2442: oled_colour = 16'b11111_111011_11011; 
		2443: oled_colour = 16'b11111_110101_10110; 
		2444: oled_colour = 16'b01100_011100_00110; 
		2445: oled_colour = 16'b01000_011011_00101; 
		2446: oled_colour = 16'b11110_110010_10100; 
		2447: oled_colour = 16'b10100_011101_01001; 
		2448: oled_colour = 16'b10100_011110_01001; 
		2449: oled_colour = 16'b11001_101011_01011; 
		2450: oled_colour = 16'b11101_101110_01100; 
		2451: oled_colour = 16'b11110_110110_00110; 
		2452: oled_colour = 16'b11101_110000_00110; 
		2453: oled_colour = 16'b11100_110000_10001; 
		2532: oled_colour = 16'b11010_101101_10110; 
		2533: oled_colour = 16'b11010_100101_01110; 
		2534: oled_colour = 16'b11110_110001_10011; 
		2535: oled_colour = 16'b11111_110111_10110; 
		2536: oled_colour = 16'b11001_101000_10010; 
		2537: oled_colour = 16'b10111_101001_10100; 
		2538: oled_colour = 16'b11111_110101_10101; 
		2539: oled_colour = 16'b11111_101111_10100; 
		2540: oled_colour = 16'b01111_011101_01000; 
		2541: oled_colour = 16'b01001_011010_00100; 
		2542: oled_colour = 16'b10101_100010_01011; 
		2543: oled_colour = 16'b10111_100001_01100; 
		2544: oled_colour = 16'b11101_101100_01111; 
		2545: oled_colour = 16'b11111_111000_00111; 
		2546: oled_colour = 16'b11110_110111_01000; 
		2547: oled_colour = 16'b11110_111010_00100; 
		2548: oled_colour = 16'b11110_111000_00101; 
		2549: oled_colour = 16'b11100_101111_01111; 
		2550: oled_colour = 16'b11111_111100_11111; 
		2627: oled_colour = 16'b11011_110011_11001; 
		2628: oled_colour = 16'b11011_101010_10000; 
		2629: oled_colour = 16'b11110_110100_10101; 
		2630: oled_colour = 16'b11011_101011_10001; 
		2631: oled_colour = 16'b11100_101111_10011; 
		2632: oled_colour = 16'b11011_101011_10000; 
		2633: oled_colour = 16'b11000_011111_01011; 
		2634: oled_colour = 16'b11101_101100_10001; 
		2635: oled_colour = 16'b11101_110000_10011; 
		2636: oled_colour = 16'b01110_100100_01100; 
		2637: oled_colour = 16'b01001_011010_00110; 
		2638: oled_colour = 16'b10101_011111_01010; 
		2639: oled_colour = 16'b11000_100011_01101; 
		2640: oled_colour = 16'b11101_101101_10100; 
		2641: oled_colour = 16'b11101_110001_01111; 
		2642: oled_colour = 16'b11101_110001_01001; 
		2643: oled_colour = 16'b11110_111001_00101; 
		2644: oled_colour = 16'b11110_110111_00101; 
		2645: oled_colour = 16'b11000_100100_01010; 
		2646: oled_colour = 16'b11101_110111_11101; 
		2723: oled_colour = 16'b11101_111000_11100; 
		2724: oled_colour = 16'b11001_101001_10001; 
		2725: oled_colour = 16'b11110_110010_10100; 
		2726: oled_colour = 16'b11110_111000_11001; 
		2727: oled_colour = 16'b11101_101111_10011; 
		2728: oled_colour = 16'b10111_100000_01100; 
		2729: oled_colour = 16'b10101_011011_01010; 
		2730: oled_colour = 16'b11011_100111_10000; 
		2731: oled_colour = 16'b11001_101000_10000; 
		2732: oled_colour = 16'b10011_101100_10000; 
		2733: oled_colour = 16'b01110_100111_01101; 
		2734: oled_colour = 16'b10001_011010_01000; 
		2735: oled_colour = 16'b10101_011101_01010; 
		2736: oled_colour = 16'b10100_011111_01010; 
		2737: oled_colour = 16'b10001_011111_01100; 
		2738: oled_colour = 16'b11011_101101_10001; 
		2739: oled_colour = 16'b11111_110111_01000; 
		2740: oled_colour = 16'b11101_110011_01010; 
		2741: oled_colour = 16'b11011_101000_01101; 
		2742: oled_colour = 16'b11001_101100_10101; 
		2819: oled_colour = 16'b11011_111000_11100; 
		2820: oled_colour = 16'b01011_011111_01001; 
		2821: oled_colour = 16'b10111_100101_01110; 
		2822: oled_colour = 16'b11010_100101_01111; 
		2823: oled_colour = 16'b11010_101010_10001; 
		2824: oled_colour = 16'b11100_101010_10000; 
		2825: oled_colour = 16'b11100_101010_10000; 
		2826: oled_colour = 16'b11110_110111_10111; 
		2827: oled_colour = 16'b11101_110011_10110; 
		2828: oled_colour = 16'b10111_100011_01110; 
		2829: oled_colour = 16'b01111_100001_01100; 
		2830: oled_colour = 16'b01010_011110_01001; 
		2831: oled_colour = 16'b01111_011110_01001; 
		2832: oled_colour = 16'b01101_011011_01001; 
		2833: oled_colour = 16'b10111_110011_11000; 
		2834: oled_colour = 16'b11111_111011_11111; 
		2835: oled_colour = 16'b11100_101011_01101; 
		2836: oled_colour = 16'b11010_100110_01101; 
		2837: oled_colour = 16'b11101_101001_10001; 
		2838: oled_colour = 16'b11001_100001_01101; 
		2839: oled_colour = 16'b11001_101010_10100; 
		2915: oled_colour = 16'b11110_111101_11110; 
		2916: oled_colour = 16'b01101_100101_01111; 
		2917: oled_colour = 16'b10100_101001_10000; 
		2918: oled_colour = 16'b11001_101010_10010; 
		2919: oled_colour = 16'b10011_101011_10001; 
		2920: oled_colour = 16'b10110_101000_01110; 
		2921: oled_colour = 16'b11101_101010_10000; 
		2922: oled_colour = 16'b11111_110001_10010; 
		2923: oled_colour = 16'b11111_110101_10110; 
		2924: oled_colour = 16'b11010_100111_01111; 
		2925: oled_colour = 16'b10101_101111_10001; 
		2926: oled_colour = 16'b11010_111100_11001; 
		2927: oled_colour = 16'b10110_110100_10101; 
		2928: oled_colour = 16'b01111_101000_10000; 
		2929: oled_colour = 16'b11101_111010_11110; 
		2931: oled_colour = 16'b11100_110100_11011; 
		2932: oled_colour = 16'b10110_100010_10000; 
		2933: oled_colour = 16'b11011_100110_01111; 
		2934: oled_colour = 16'b11111_110011_10101; 
		2935: oled_colour = 16'b11011_101100_10001; 
		2936: oled_colour = 16'b11010_101101_10110; 
		3013: oled_colour = 16'b10110_101101_10101; 
		3014: oled_colour = 16'b10011_100110_01111; 
		3015: oled_colour = 16'b10000_101010_10000; 
		3016: oled_colour = 16'b10000_101111_10000; 
		3017: oled_colour = 16'b10111_110011_10011; 
		3018: oled_colour = 16'b11001_101101_10000; 
		3019: oled_colour = 16'b11101_101011_10001; 
		3020: oled_colour = 16'b10100_101000_01111; 
		3021: oled_colour = 16'b01101_100011_01011; 
		3022: oled_colour = 16'b11010_110010_10010; 
		3023: oled_colour = 16'b11111_111010_11000; 
		3024: oled_colour = 16'b11010_110000_10010; 
		3025: oled_colour = 16'b10100_100010_01110; 
		3026: oled_colour = 16'b11111_111101_11111; 
		3028: oled_colour = 16'b11111_111110_11111; 
		3029: oled_colour = 16'b11001_101011_10100; 
		3030: oled_colour = 16'b11100_101100_10000; 
		3031: oled_colour = 16'b11111_110111_10101; 
		3032: oled_colour = 16'b11010_101010_10001; 
		3033: oled_colour = 16'b11101_111000_11100; 
		3110: oled_colour = 16'b11001_110101_11010; 
		3111: oled_colour = 16'b01111_100100_01110; 
		3112: oled_colour = 16'b00111_011011_01000; 
		3113: oled_colour = 16'b01100_100001_01011; 
		3114: oled_colour = 16'b10000_100110_01011; 
		3115: oled_colour = 16'b11011_111011_10111; 
		3116: oled_colour = 16'b11110_111110_11100; 
		3117: oled_colour = 16'b10011_100010_01100; 
		3118: oled_colour = 16'b10100_011000_01001; 
		3119: oled_colour = 16'b11001_101011_10000; 
		3120: oled_colour = 16'b11111_110111_10100; 
		3121: oled_colour = 16'b11001_110001_10011; 
		3122: oled_colour = 16'b10001_101001_10001; 
		3123: oled_colour = 16'b11111_111101_11111; 
		3126: oled_colour = 16'b11010_101110_10111; 
		3127: oled_colour = 16'b11010_100110_01111; 
		3128: oled_colour = 16'b11101_101101_10000; 
		3129: oled_colour = 16'b11010_101011_10100; 
		3208: oled_colour = 16'b11100_111010_11100; 
		3209: oled_colour = 16'b01110_011011_01010; 
		3210: oled_colour = 16'b10001_011101_01001; 
		3211: oled_colour = 16'b11101_101110_10010; 
		3212: oled_colour = 16'b11111_110100_10100; 
		3213: oled_colour = 16'b11110_110000_10010; 
		3214: oled_colour = 16'b01101_011110_01001; 
		3215: oled_colour = 16'b01100_100011_01100; 
		3216: oled_colour = 16'b10110_110110_10011; 
		3217: oled_colour = 16'b11110_111111_11011; 
		3218: oled_colour = 16'b10010_101111_10000; 
		3219: oled_colour = 16'b10000_101000_10010; 
		3223: oled_colour = 16'b11011_110010_11010; 
		3224: oled_colour = 16'b11011_101001_10000; 
		3225: oled_colour = 16'b11110_110011_10100; 
		3226: oled_colour = 16'b11011_110000_10110; 
		3305: oled_colour = 16'b11011_110111_11011; 
		3306: oled_colour = 16'b01011_011000_00111; 
		3307: oled_colour = 16'b11001_101111_10110; 
		3308: oled_colour = 16'b11100_110110_11001; 
		3309: oled_colour = 16'b10111_110101_10101; 
		3310: oled_colour = 16'b01110_101011_01111; 
		3311: oled_colour = 16'b01000_010110_00100; 
		3312: oled_colour = 16'b01011_010100_00011; 
		3313: oled_colour = 16'b01101_011110_01000; 
		3314: oled_colour = 16'b10000_100010_01011; 
		3315: oled_colour = 16'b10000_011100_01010; 
		3316: oled_colour = 16'b11111_111110_11111; 
		3319: oled_colour = 16'b11111_111101_11111; 
		3320: oled_colour = 16'b11001_101001_10011; 
		3321: oled_colour = 16'b11100_110000_10101; 
		3322: oled_colour = 16'b11001_100110_10000; 
		3323: oled_colour = 16'b11000_101001_10011; 
		3402: oled_colour = 16'b10110_101111_10110; 
		3403: oled_colour = 16'b01011_010101_00100; 
		3404: oled_colour = 16'b01011_010100_00011; 
		3405: oled_colour = 16'b10010_100010_01011; 
		3406: oled_colour = 16'b10011_011111_01011; 
		3407: oled_colour = 16'b01101_011001_01000; 
		3408: oled_colour = 16'b01100_100000_01100; 
		3409: oled_colour = 16'b01100_011001_00111; 
		3410: oled_colour = 16'b11000_011110_01011; 
		3411: oled_colour = 16'b10001_010101_00110; 
		3412: oled_colour = 16'b10011_011111_01101; 
		3416: oled_colour = 16'b11010_101111_10111; 
		3417: oled_colour = 16'b11111_111101_11111; 
		3418: oled_colour = 16'b11111_111110_11111; 
		3419: oled_colour = 16'b11010_110000_10111; 
		3420: oled_colour = 16'b11101_110111_11100; 
		3499: oled_colour = 16'b11000_110000_10110; 
		3500: oled_colour = 16'b01101_011011_01001; 
		3501: oled_colour = 16'b10111_011110_01011; 
		3502: oled_colour = 16'b10011_011001_00110; 
		3503: oled_colour = 16'b10001_011000_01000; 
		3505: oled_colour = 16'b11011_110000_11000; 
		3506: oled_colour = 16'b10011_011001_01001; 
		3507: oled_colour = 16'b11000_100011_01100; 
		3508: oled_colour = 16'b01111_010011_00100; 
		3509: oled_colour = 16'b10010_011101_01011; 
		3510: oled_colour = 16'b10111_101001_10011; 
		3511: oled_colour = 16'b11011_101101_10101; 
		3512: oled_colour = 16'b11100_110000_10111; 
		3513: oled_colour = 16'b11101_110111_11011; 
		3596: oled_colour = 16'b11111_111011_11110; 
		3597: oled_colour = 16'b01111_010110_00111; 
		3598: oled_colour = 16'b01010_001110_00001; 
		3599: oled_colour = 16'b01101_010011_00011; 
		3600: oled_colour = 16'b10001_011011_01001; 
		3601: oled_colour = 16'b10100_011111_01101; 
		3602: oled_colour = 16'b11000_100000_01100; 
		3603: oled_colour = 16'b11100_100101_01111; 
		3604: oled_colour = 16'b10010_011010_01000; 
		3605: oled_colour = 16'b01011_001110_00001; 
		3606: oled_colour = 16'b01110_010000_00010; 
		3607: oled_colour = 16'b10101_011001_01001; 
		3608: oled_colour = 16'b10101_011001_01000; 
		3609: oled_colour = 16'b10011_011001_01010; 
		3610: oled_colour = 16'b11101_111001_11101; 
		3693: oled_colour = 16'b11100_110111_11011; 
		3694: oled_colour = 16'b01101_010100_00100; 
		3695: oled_colour = 16'b01100_010000_00001; 
		3696: oled_colour = 16'b01011_001111_00001; 
		3697: oled_colour = 16'b01101_010000_00001; 
		3698: oled_colour = 16'b10001_011000_01000; 
		3699: oled_colour = 16'b10110_100010_01111; 
		3700: oled_colour = 16'b10100_011010_01001; 
		3701: oled_colour = 16'b10100_011100_01010; 
		3702: oled_colour = 16'b10010_011110_01011; 
		3703: oled_colour = 16'b10110_100011_01111; 
		3704: oled_colour = 16'b11001_101100_10101; 
		3705: oled_colour = 16'b11100_110101_11011; 
		3790: oled_colour = 16'b11011_110011_11001; 
		3791: oled_colour = 16'b10110_011111_01011; 
		3792: oled_colour = 16'b10101_011011_01001; 
		3793: oled_colour = 16'b10010_011010_01001; 
		3794: oled_colour = 16'b11100_110111_11011; 
		3796: oled_colour = 16'b11100_110011_11010; 
		3797: oled_colour = 16'b11101_110111_11100; 
		3887: oled_colour = 16'b11001_101100_10101; 
		3888: oled_colour = 16'b10101_011100_01010; 
		3889: oled_colour = 16'b11010_101100_10101; 
		3984: oled_colour = 16'b11111_111101_11111; 
		default: oled_colour = 16'b00000_000000_00000; 
	endcase
end

endmodule