module Gui_State1(
    input [12:0] pixel_index, 
    output reg [15:0] oled_colour 
); 

always@(pixel_index) 
begin
	case(pixel_index)
		1872: oled_colour = 16'b11110_111001_11100; 
		1873: oled_colour = 16'b11110_111000_11010; 
		1874: oled_colour = 16'b11111_111100_11100; 
		1875: oled_colour = 16'b11111_111101_11001; 
		1876: oled_colour = 16'b11111_111110_11001; 
		1877: oled_colour = 16'b11111_111101_11010; 
		1878: oled_colour = 16'b11111_111101_11011; 
		1879: oled_colour = 16'b11111_111110_11101; 
		1880: oled_colour = 16'b11111_111110_11101; 
		1881: oled_colour = 16'b11111_111110_11111; 
		1965: oled_colour = 16'b11111_111110_11111; 
		1966: oled_colour = 16'b11111_111101_11110; 
		1969: oled_colour = 16'b11110_110100_10101; 
		1970: oled_colour = 16'b11101_101110_01011; 
		1971: oled_colour = 16'b11110_110101_01010; 
		1972: oled_colour = 16'b11101_110100_00101; 
		1973: oled_colour = 16'b11110_110100_01010; 
		1974: oled_colour = 16'b11110_110010_00111; 
		1975: oled_colour = 16'b11110_110100_01101; 
		1976: oled_colour = 16'b11111_111001_11000; 
		1977: oled_colour = 16'b11111_111100_11110; 
		2060: oled_colour = 16'b11101_110101_11010; 
		2061: oled_colour = 16'b11011_101101_10011; 
		2062: oled_colour = 16'b11101_110011_11000; 
		2063: oled_colour = 16'b11011_110001_10101; 
		2064: oled_colour = 16'b10111_110000_10101; 
		2065: oled_colour = 16'b11001_101011_10100; 
		2066: oled_colour = 16'b11010_100111_01100; 
		2067: oled_colour = 16'b11101_110000_01100; 
		2068: oled_colour = 16'b11100_101111_10010; 
		2069: oled_colour = 16'b11101_110001_01111; 
		2070: oled_colour = 16'b11101_110010_10011; 
		2155: oled_colour = 16'b11111_111101_11110; 
		2156: oled_colour = 16'b11010_101010_10010; 
		2157: oled_colour = 16'b11101_101111_10011; 
		2158: oled_colour = 16'b11101_110011_10110; 
		2159: oled_colour = 16'b11100_101011_10000; 
		2160: oled_colour = 16'b01110_100001_01001; 
		2161: oled_colour = 16'b01110_010111_00101; 
		2162: oled_colour = 16'b11001_100110_10000; 
		2163: oled_colour = 16'b11010_100111_01110; 
		2164: oled_colour = 16'b11011_101100_10100; 
		2165: oled_colour = 16'b11001_101001_10011; 
		2166: oled_colour = 16'b11011_101100_10011; 
		2167: oled_colour = 16'b11111_111110_11111; 
		2168: oled_colour = 16'b11111_111100_11110; 
		2169: oled_colour = 16'b11011_110000_10111; 
		2170: oled_colour = 16'b11110_111001_11100; 
		2251: oled_colour = 16'b11101_111011_11101; 
		2252: oled_colour = 16'b10110_100001_01100; 
		2253: oled_colour = 16'b10111_011101_01011; 
		2254: oled_colour = 16'b10111_100100_10001; 
		2255: oled_colour = 16'b11011_101001_10001; 
		2256: oled_colour = 16'b10011_011101_01011; 
		2257: oled_colour = 16'b10110_011111_01011; 
		2258: oled_colour = 16'b11111_101101_10011; 
		2259: oled_colour = 16'b11001_100110_01111; 
		2260: oled_colour = 16'b11011_101100_10011; 
		2261: oled_colour = 16'b11000_101010_10001; 
		2262: oled_colour = 16'b11011_101100_10001; 
		2263: oled_colour = 16'b11110_110101_11010; 
		2264: oled_colour = 16'b11010_101111_10110; 
		2265: oled_colour = 16'b10110_100001_01100; 
		2266: oled_colour = 16'b10111_100010_01110; 
		2267: oled_colour = 16'b11110_110111_11011; 
		2347: oled_colour = 16'b11011_111010_11100; 
		2348: oled_colour = 16'b01111_011100_00111; 
		2349: oled_colour = 16'b11101_100111_01111; 
		2350: oled_colour = 16'b11100_101100_10010; 
		2351: oled_colour = 16'b11001_101000_10000; 
		2352: oled_colour = 16'b11000_100100_01101; 
		2353: oled_colour = 16'b11110_101110_10010; 
		2354: oled_colour = 16'b11001_100110_01111; 
		2355: oled_colour = 16'b10100_011101_01010; 
		2356: oled_colour = 16'b10101_100000_01100; 
		2357: oled_colour = 16'b10011_100000_01011; 
		2358: oled_colour = 16'b11011_101100_10011; 
		2359: oled_colour = 16'b11001_101000_10001; 
		2360: oled_colour = 16'b11000_100011_01110; 
		2361: oled_colour = 16'b11001_100111_01111; 
		2362: oled_colour = 16'b10111_100010_01101; 
		2363: oled_colour = 16'b11100_110101_11010; 
		2443: oled_colour = 16'b11111_111110_11111; 
		2444: oled_colour = 16'b01101_011101_01001; 
		2445: oled_colour = 16'b11000_100001_01101; 
		2446: oled_colour = 16'b11001_100111_01111; 
		2447: oled_colour = 16'b11101_110101_10111; 
		2448: oled_colour = 16'b11111_111001_11000; 
		2449: oled_colour = 16'b11000_100110_01101; 
		2450: oled_colour = 16'b01100_011011_01000; 
		2451: oled_colour = 16'b10000_011110_01001; 
		2452: oled_colour = 16'b01101_011111_01001; 
		2453: oled_colour = 16'b01001_011001_00110; 
		2454: oled_colour = 16'b11001_100111_10001; 
		2455: oled_colour = 16'b11011_100110_01111; 
		2456: oled_colour = 16'b11100_101010_10000; 
		2457: oled_colour = 16'b11001_101001_10010; 
		2458: oled_colour = 16'b11111_111100_11110; 
		2540: oled_colour = 16'b01110_100100_01101; 
		2541: oled_colour = 16'b10011_011011_01000; 
		2542: oled_colour = 16'b11111_110101_10111; 
		2543: oled_colour = 16'b11101_101111_10101; 
		2544: oled_colour = 16'b10111_011111_01011; 
		2545: oled_colour = 16'b01001_011000_00101; 
		2546: oled_colour = 16'b01000_011110_01000; 
		2547: oled_colour = 16'b00111_011011_00110; 
		2548: oled_colour = 16'b01110_100100_01101; 
		2549: oled_colour = 16'b10000_011000_00111; 
		2550: oled_colour = 16'b11010_100100_01110; 
		2551: oled_colour = 16'b11111_110110_10111; 
		2552: oled_colour = 16'b11011_101011_10001; 
		2553: oled_colour = 16'b11111_111100_11110; 
		2636: oled_colour = 16'b10011_101010_10001; 
		2637: oled_colour = 16'b01110_011010_00111; 
		2638: oled_colour = 16'b11000_100110_01110; 
		2639: oled_colour = 16'b01010_010101_00011; 
		2640: oled_colour = 16'b00100_010100_00001; 
		2641: oled_colour = 16'b00001_010011_00001; 
		2642: oled_colour = 16'b00001_010011_00001; 
		2643: oled_colour = 16'b10100_101101_10011; 
		2645: oled_colour = 16'b11011_101101_10101; 
		2646: oled_colour = 16'b11011_101100_10011; 
		2647: oled_colour = 16'b11010_101001_10001; 
		2648: oled_colour = 16'b11100_110100_11001; 
		2732: oled_colour = 16'b10011_100111_10000; 
		2733: oled_colour = 16'b01100_010111_00110; 
		2734: oled_colour = 16'b01110_011000_00110; 
		2735: oled_colour = 16'b01011_011010_00101; 
		2736: oled_colour = 16'b01011_011010_00101; 
		2737: oled_colour = 16'b01100_100000_01001; 
		2738: oled_colour = 16'b01010_010110_00100; 
		2739: oled_colour = 16'b11101_111000_11100; 
		2742: oled_colour = 16'b11111_111011_11101; 
		2743: oled_colour = 16'b11111_111100_11110; 
		2827: oled_colour = 16'b11101_111001_11101; 
		2828: oled_colour = 16'b10011_011011_01001; 
		2829: oled_colour = 16'b10001_100100_01101; 
		2830: oled_colour = 16'b10001_011001_01000; 
		2831: oled_colour = 16'b10011_011000_01000; 
		2832: oled_colour = 16'b01110_011111_01010; 
		2833: oled_colour = 16'b01010_011101_01000; 
		2834: oled_colour = 16'b01111_010110_00101; 
		2835: oled_colour = 16'b11101_110111_11010; 
		2923: oled_colour = 16'b11011_110100_11000; 
		2924: oled_colour = 16'b10010_100100_01110; 
		2925: oled_colour = 16'b10111_110000_10010; 
		2926: oled_colour = 16'b10110_101010_10000; 
		2927: oled_colour = 16'b10001_011001_01000; 
		2928: oled_colour = 16'b01001_011000_00101; 
		2929: oled_colour = 16'b00101_011000_00100; 
		2930: oled_colour = 16'b01010_010100_00011; 
		2931: oled_colour = 16'b10111_110001_10110; 
		3019: oled_colour = 16'b11101_111100_11100; 
		3020: oled_colour = 16'b10011_101111_10011; 
		3021: oled_colour = 16'b10011_110011_10010; 
		3022: oled_colour = 16'b11010_111101_10100; 
		3023: oled_colour = 16'b10001_101100_01111; 
		3024: oled_colour = 16'b01000_011000_00100; 
		3025: oled_colour = 16'b00110_011001_00100; 
		3026: oled_colour = 16'b01010_011001_00110; 
		3027: oled_colour = 16'b10101_110000_10110; 
		3115: oled_colour = 16'b11101_111101_11101; 
		3116: oled_colour = 16'b10111_110001_10100; 
		3117: oled_colour = 16'b11001_101111_10011; 
		3118: oled_colour = 16'b11110_110111_10111; 
		3119: oled_colour = 16'b11001_110010_10110; 
		3120: oled_colour = 16'b10000_100111_01111; 
		3121: oled_colour = 16'b00101_010100_00010; 
		3122: oled_colour = 16'b10000_100001_01010; 
		3123: oled_colour = 16'b11010_110001_10101; 
		3211: oled_colour = 16'b11101_110111_11011; 
		3212: oled_colour = 16'b11100_101111_10100; 
		3213: oled_colour = 16'b11100_110000_10101; 
		3214: oled_colour = 16'b11101_101011_10010; 
		3215: oled_colour = 16'b11111_110100_10011; 
		3216: oled_colour = 16'b11001_101110_10010; 
		3217: oled_colour = 16'b00101_010110_00100; 
		3218: oled_colour = 16'b10111_101001_10001; 
		3219: oled_colour = 16'b11110_110101_11000; 
		3220: oled_colour = 16'b11110_111010_11101; 
		3307: oled_colour = 16'b11110_111001_11100; 
		3308: oled_colour = 16'b10010_101010_10001; 
		3309: oled_colour = 16'b10010_101111_10010; 
		3310: oled_colour = 16'b11011_110011_10010; 
		3311: oled_colour = 16'b11110_110100_10010; 
		3312: oled_colour = 16'b10110_110110_10010; 
		3313: oled_colour = 16'b01001_011100_01000; 
		3314: oled_colour = 16'b10110_110001_10010; 
		3315: oled_colour = 16'b11011_110101_10010; 
		3316: oled_colour = 16'b11100_101111_10101; 
		3404: oled_colour = 16'b11001_110110_11010; 
		3405: oled_colour = 16'b01100_100011_01011; 
		3406: oled_colour = 16'b10011_101011_01101; 
		3407: oled_colour = 16'b11100_110001_10011; 
		3408: oled_colour = 16'b11100_110100_10101; 
		3409: oled_colour = 16'b01100_100000_01011; 
		3410: oled_colour = 16'b10100_101101_10000; 
		3411: oled_colour = 16'b11111_111001_10111; 
		3412: oled_colour = 16'b11011_101111_10011; 
		3413: oled_colour = 16'b11111_111100_11110; 
		3501: oled_colour = 16'b10101_100100_01110; 
		3502: oled_colour = 16'b01100_011010_00111; 
		3503: oled_colour = 16'b10111_110011_10011; 
		3504: oled_colour = 16'b11000_111010_10110; 
		3505: oled_colour = 16'b01000_011101_01000; 
		3506: oled_colour = 16'b10000_101100_01110; 
		3507: oled_colour = 16'b11110_111100_11010; 
		3508: oled_colour = 16'b10100_100100_01101; 
		3509: oled_colour = 16'b11101_111000_11011; 
		3596: oled_colour = 16'b11110_111100_11110; 
		3597: oled_colour = 16'b10110_100111_01110; 
		3598: oled_colour = 16'b11000_101101_10010; 
		3599: oled_colour = 16'b10101_110011_10101; 
		3600: oled_colour = 16'b10111_110010_10011; 
		3601: oled_colour = 16'b10000_011010_01000; 
		3602: oled_colour = 16'b01111_100111_10000; 
		3603: oled_colour = 16'b10011_101110_10000; 
		3604: oled_colour = 16'b10110_101011_10010; 
		3605: oled_colour = 16'b11111_111110_11111; 
		3692: oled_colour = 16'b11111_111100_11110; 
		3693: oled_colour = 16'b01110_011110_01001; 
		3694: oled_colour = 16'b10100_110001_10011; 
		3695: oled_colour = 16'b11001_110000_10100; 
		3696: oled_colour = 16'b10001_100000_01011; 
		3697: oled_colour = 16'b01011_010110_00101; 
		3698: oled_colour = 16'b10001_100000_01011; 
		3699: oled_colour = 16'b11010_110011_10111; 
		3789: oled_colour = 16'b10101_101001_10001; 
		3790: oled_colour = 16'b01010_010110_00100; 
		3791: oled_colour = 16'b01011_011101_00111; 
		3792: oled_colour = 16'b01010_010011_00010; 
		3793: oled_colour = 16'b01111_010110_00101; 
		3794: oled_colour = 16'b10110_101010_10010; 
		3885: oled_colour = 16'b10111_101011_10011; 
		3886: oled_colour = 16'b10001_010110_00101; 
		3887: oled_colour = 16'b10001_010110_00101; 
		3888: oled_colour = 16'b01110_010001_00010; 
		3889: oled_colour = 16'b10110_100000_01100; 
		3981: oled_colour = 16'b10111_101010_10010; 
		3982: oled_colour = 16'b10001_010110_00101; 
		3983: oled_colour = 16'b01111_010101_00100; 
		3984: oled_colour = 16'b01101_010001_00010; 
		3985: oled_colour = 16'b10100_011101_01010; 
		3986: oled_colour = 16'b11111_111110_11111; 
		4077: oled_colour = 16'b10111_101011_10011; 
		4078: oled_colour = 16'b10010_011000_00110; 
		4079: oled_colour = 16'b01111_010100_00100; 
		4080: oled_colour = 16'b10100_011101_01001; 
		4081: oled_colour = 16'b11010_100111_01111; 
		4082: oled_colour = 16'b11100_110011_11000; 
		4173: oled_colour = 16'b11011_110001_10111; 
		4174: oled_colour = 16'b11001_100010_01100; 
		4175: oled_colour = 16'b11001_100100_01110; 
		4176: oled_colour = 16'b11011_101100_10100; 
		4177: oled_colour = 16'b11100_101111_10100; 
		4178: oled_colour = 16'b11111_111001_11100; 
		4270: oled_colour = 16'b11101_110110_11010; 
		4271: oled_colour = 16'b11111_111010_11100; 
		default: oled_colour = 16'b00000_000000_00000; 
	endcase
end

endmodule