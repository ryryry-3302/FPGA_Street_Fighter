module Gui_b2(
    input [12:0] pixel_index, 
    output reg [15:0] oled_colour 
); 

always@(pixel_index) 
begin
	case(pixel_index)
		0: oled_colour = 16'b00001_000001_00001; 
		1: oled_colour = 16'b00001_000001_00001; 
		2: oled_colour = 16'b00001_000001_00001; 
		3: oled_colour = 16'b00001_000001_00001; 
		4: oled_colour = 16'b00001_000001_00001; 
		5: oled_colour = 16'b00001_000001_00001; 
		6: oled_colour = 16'b00001_000001_00001; 
		7: oled_colour = 16'b00001_000001_00001; 
		8: oled_colour = 16'b00001_000001_00001; 
		9: oled_colour = 16'b00001_000001_00001; 
		10: oled_colour = 16'b00001_000001_00001; 
		11: oled_colour = 16'b00001_000001_00001; 
		12: oled_colour = 16'b00001_000001_00001; 
		13: oled_colour = 16'b00001_000001_00001; 
		14: oled_colour = 16'b00001_000001_00001; 
		15: oled_colour = 16'b00001_000001_00001; 
		16: oled_colour = 16'b00001_000001_00001; 
		17: oled_colour = 16'b00001_000001_00001; 
		18: oled_colour = 16'b00001_000001_00001; 
		19: oled_colour = 16'b00001_000001_00001; 
		20: oled_colour = 16'b00001_000001_00001; 
		21: oled_colour = 16'b00001_000001_00001; 
		22: oled_colour = 16'b00001_000001_00001; 
		23: oled_colour = 16'b00001_000001_00001; 
		24: oled_colour = 16'b00001_000001_00001; 
		25: oled_colour = 16'b00001_000001_00001; 
		26: oled_colour = 16'b00001_000001_00001; 
		27: oled_colour = 16'b00001_000001_00001; 
		28: oled_colour = 16'b00001_000001_00001; 
		29: oled_colour = 16'b00001_000001_00001; 
		30: oled_colour = 16'b00001_000001_00001; 
		31: oled_colour = 16'b00001_000001_00001; 
		32: oled_colour = 16'b00001_000001_00001; 
		33: oled_colour = 16'b00001_000001_00001; 
		34: oled_colour = 16'b00001_000001_00001; 
		35: oled_colour = 16'b00001_000001_00001; 
		36: oled_colour = 16'b00001_000001_00001; 
		37: oled_colour = 16'b00001_000001_00001; 
		38: oled_colour = 16'b00001_000001_00001; 
		39: oled_colour = 16'b00001_000001_00001; 
		40: oled_colour = 16'b00001_000001_00001; 
		41: oled_colour = 16'b00001_000001_00001; 
		42: oled_colour = 16'b00001_000001_00001; 
		43: oled_colour = 16'b00001_000001_00001; 
		44: oled_colour = 16'b00001_000001_00001; 
		45: oled_colour = 16'b00001_000001_00001; 
		46: oled_colour = 16'b00001_000001_00001; 
		47: oled_colour = 16'b00001_000001_00001; 
		48: oled_colour = 16'b00001_000001_00001; 
		49: oled_colour = 16'b00001_000001_00001; 
		50: oled_colour = 16'b00001_000001_00001; 
		51: oled_colour = 16'b00001_000001_00001; 
		52: oled_colour = 16'b00001_000001_00001; 
		53: oled_colour = 16'b00001_000001_00001; 
		54: oled_colour = 16'b00001_000001_00001; 
		55: oled_colour = 16'b00001_000001_00001; 
		56: oled_colour = 16'b00001_000001_00001; 
		57: oled_colour = 16'b00001_000001_00001; 
		58: oled_colour = 16'b00001_000001_00001; 
		59: oled_colour = 16'b00001_000001_00001; 
		60: oled_colour = 16'b00001_000001_00001; 
		61: oled_colour = 16'b00001_000001_00001; 
		62: oled_colour = 16'b00001_000001_00001; 
		63: oled_colour = 16'b00001_000001_00001; 
		64: oled_colour = 16'b00001_000001_00001; 
		65: oled_colour = 16'b00001_000001_00001; 
		66: oled_colour = 16'b00001_000001_00001; 
		67: oled_colour = 16'b00001_000001_00001; 
		68: oled_colour = 16'b00001_000001_00001; 
		69: oled_colour = 16'b00001_000001_00001; 
		70: oled_colour = 16'b00001_000001_00001; 
		71: oled_colour = 16'b00001_000001_00001; 
		72: oled_colour = 16'b00001_000001_00001; 
		73: oled_colour = 16'b00001_000001_00001; 
		74: oled_colour = 16'b00001_000001_00001; 
		75: oled_colour = 16'b00001_000001_00001; 
		76: oled_colour = 16'b00001_000001_00001; 
		77: oled_colour = 16'b00001_000001_00001; 
		78: oled_colour = 16'b00001_000001_00001; 
		79: oled_colour = 16'b00001_000001_00001; 
		80: oled_colour = 16'b00001_000001_00001; 
		81: oled_colour = 16'b00001_000001_00001; 
		82: oled_colour = 16'b00001_000001_00001; 
		83: oled_colour = 16'b00001_000001_00001; 
		84: oled_colour = 16'b00001_000001_00001; 
		85: oled_colour = 16'b00001_000001_00001; 
		86: oled_colour = 16'b00001_000001_00001; 
		87: oled_colour = 16'b00001_000001_00001; 
		88: oled_colour = 16'b00001_000001_00001; 
		89: oled_colour = 16'b00001_000001_00001; 
		90: oled_colour = 16'b00001_000001_00001; 
		91: oled_colour = 16'b00001_000001_00001; 
		92: oled_colour = 16'b00001_000001_00001; 
		93: oled_colour = 16'b00001_000001_00001; 
		94: oled_colour = 16'b00001_000001_00001; 
		95: oled_colour = 16'b00001_000001_00001; 
		96: oled_colour = 16'b00001_000001_00001; 
		97: oled_colour = 16'b00001_000001_00001; 
		98: oled_colour = 16'b00001_000001_00001; 
		99: oled_colour = 16'b00001_000001_00001; 
		100: oled_colour = 16'b00001_000001_00001; 
		101: oled_colour = 16'b00001_000001_00001; 
		102: oled_colour = 16'b00001_000001_00001; 
		103: oled_colour = 16'b00001_000001_00001; 
		104: oled_colour = 16'b00001_000001_00001; 
		105: oled_colour = 16'b00001_000001_00001; 
		106: oled_colour = 16'b00001_000001_00001; 
		107: oled_colour = 16'b00001_000001_00001; 
		108: oled_colour = 16'b00001_000001_00001; 
		109: oled_colour = 16'b00001_000001_00001; 
		110: oled_colour = 16'b00001_000001_00001; 
		111: oled_colour = 16'b00001_000001_00001; 
		112: oled_colour = 16'b00001_000001_00001; 
		113: oled_colour = 16'b00001_000001_00001; 
		114: oled_colour = 16'b00001_000001_00001; 
		115: oled_colour = 16'b00001_000001_00001; 
		116: oled_colour = 16'b00001_000001_00001; 
		117: oled_colour = 16'b00001_000001_00001; 
		118: oled_colour = 16'b00001_000001_00001; 
		119: oled_colour = 16'b00001_000001_00001; 
		120: oled_colour = 16'b00001_000001_00001; 
		121: oled_colour = 16'b00001_000001_00001; 
		122: oled_colour = 16'b00001_000001_00001; 
		123: oled_colour = 16'b00001_000001_00001; 
		124: oled_colour = 16'b00001_000001_00001; 
		125: oled_colour = 16'b00001_000001_00001; 
		126: oled_colour = 16'b00001_000001_00001; 
		127: oled_colour = 16'b00001_000001_00001; 
		128: oled_colour = 16'b00001_000001_00001; 
		129: oled_colour = 16'b00001_000001_00001; 
		130: oled_colour = 16'b00001_000001_00001; 
		131: oled_colour = 16'b00001_000001_00001; 
		132: oled_colour = 16'b00001_000001_00001; 
		133: oled_colour = 16'b00001_000001_00001; 
		134: oled_colour = 16'b00001_000001_00001; 
		135: oled_colour = 16'b00001_000001_00001; 
		136: oled_colour = 16'b00001_000001_00001; 
		137: oled_colour = 16'b00001_000001_00001; 
		138: oled_colour = 16'b00001_000001_00001; 
		139: oled_colour = 16'b00001_000001_00001; 
		140: oled_colour = 16'b00001_000001_00001; 
		141: oled_colour = 16'b00001_000001_00001; 
		142: oled_colour = 16'b00001_000001_00001; 
		143: oled_colour = 16'b00001_000001_00001; 
		144: oled_colour = 16'b00001_000001_00001; 
		145: oled_colour = 16'b00001_000001_00001; 
		146: oled_colour = 16'b00001_000001_00001; 
		147: oled_colour = 16'b00001_000001_00001; 
		148: oled_colour = 16'b00001_000001_00001; 
		149: oled_colour = 16'b00001_000001_00001; 
		150: oled_colour = 16'b00001_000001_00001; 
		151: oled_colour = 16'b00001_000001_00001; 
		152: oled_colour = 16'b00001_000001_00001; 
		153: oled_colour = 16'b00001_000001_00001; 
		154: oled_colour = 16'b00001_000001_00001; 
		155: oled_colour = 16'b00001_000001_00001; 
		156: oled_colour = 16'b00001_000001_00001; 
		157: oled_colour = 16'b00001_000001_00001; 
		158: oled_colour = 16'b00001_000001_00001; 
		159: oled_colour = 16'b00001_000001_00001; 
		160: oled_colour = 16'b00001_000001_00001; 
		161: oled_colour = 16'b00001_000001_00001; 
		162: oled_colour = 16'b00001_000001_00001; 
		163: oled_colour = 16'b00001_000001_00001; 
		164: oled_colour = 16'b00001_000001_00001; 
		165: oled_colour = 16'b00001_000001_00001; 
		166: oled_colour = 16'b00001_000001_00001; 
		167: oled_colour = 16'b00001_000001_00001; 
		168: oled_colour = 16'b00001_000001_00001; 
		169: oled_colour = 16'b00001_000001_00001; 
		170: oled_colour = 16'b00001_000001_00001; 
		171: oled_colour = 16'b00001_000001_00001; 
		172: oled_colour = 16'b00001_000001_00001; 
		173: oled_colour = 16'b00001_000001_00001; 
		174: oled_colour = 16'b00001_000001_00001; 
		175: oled_colour = 16'b00001_000001_00001; 
		176: oled_colour = 16'b00001_000001_00001; 
		177: oled_colour = 16'b00001_000001_00001; 
		178: oled_colour = 16'b00001_000001_00001; 
		179: oled_colour = 16'b00001_000001_00001; 
		180: oled_colour = 16'b00001_000001_00001; 
		181: oled_colour = 16'b00001_000001_00001; 
		182: oled_colour = 16'b00001_000001_00001; 
		183: oled_colour = 16'b00001_000001_00001; 
		184: oled_colour = 16'b00001_000001_00001; 
		185: oled_colour = 16'b00001_000001_00001; 
		186: oled_colour = 16'b00001_000001_00001; 
		187: oled_colour = 16'b00001_000001_00001; 
		188: oled_colour = 16'b00001_000001_00001; 
		189: oled_colour = 16'b00001_000001_00001; 
		190: oled_colour = 16'b00001_000001_00001; 
		191: oled_colour = 16'b00001_000001_00001; 
		192: oled_colour = 16'b00001_000001_00001; 
		193: oled_colour = 16'b00001_000001_00001; 
		194: oled_colour = 16'b00001_000001_00001; 
		195: oled_colour = 16'b00001_000001_00001; 
		196: oled_colour = 16'b00001_000001_00001; 
		197: oled_colour = 16'b00001_000001_00001; 
		198: oled_colour = 16'b00001_000001_00001; 
		199: oled_colour = 16'b00001_000001_00001; 
		200: oled_colour = 16'b00001_000001_00001; 
		201: oled_colour = 16'b00001_000001_00001; 
		202: oled_colour = 16'b00001_000001_00001; 
		203: oled_colour = 16'b00001_000001_00001; 
		204: oled_colour = 16'b00001_000001_00001; 
		205: oled_colour = 16'b00001_000001_00001; 
		206: oled_colour = 16'b00001_000001_00001; 
		207: oled_colour = 16'b00001_000001_00001; 
		208: oled_colour = 16'b00001_000001_00001; 
		209: oled_colour = 16'b00001_000001_00001; 
		210: oled_colour = 16'b00001_000001_00001; 
		211: oled_colour = 16'b00001_000001_00001; 
		212: oled_colour = 16'b00001_000001_00001; 
		213: oled_colour = 16'b00001_000001_00001; 
		214: oled_colour = 16'b00001_000001_00001; 
		215: oled_colour = 16'b00001_000001_00001; 
		216: oled_colour = 16'b00001_000001_00001; 
		217: oled_colour = 16'b00001_000001_00001; 
		218: oled_colour = 16'b00001_000001_00001; 
		219: oled_colour = 16'b00001_000001_00001; 
		220: oled_colour = 16'b00001_000001_00001; 
		221: oled_colour = 16'b00001_000001_00001; 
		222: oled_colour = 16'b00001_000001_00001; 
		223: oled_colour = 16'b00001_000001_00001; 
		224: oled_colour = 16'b00001_000001_00001; 
		225: oled_colour = 16'b00001_000001_00001; 
		226: oled_colour = 16'b00001_000001_00001; 
		227: oled_colour = 16'b00001_000001_00001; 
		228: oled_colour = 16'b00001_000001_00001; 
		229: oled_colour = 16'b00001_000001_00001; 
		230: oled_colour = 16'b00001_000001_00001; 
		231: oled_colour = 16'b00001_000001_00001; 
		232: oled_colour = 16'b00001_000001_00001; 
		233: oled_colour = 16'b00001_000001_00001; 
		234: oled_colour = 16'b00001_000001_00001; 
		235: oled_colour = 16'b00001_000001_00001; 
		236: oled_colour = 16'b00001_000001_00001; 
		237: oled_colour = 16'b00001_000001_00001; 
		238: oled_colour = 16'b00001_000001_00001; 
		239: oled_colour = 16'b00001_000001_00001; 
		240: oled_colour = 16'b00001_000001_00001; 
		241: oled_colour = 16'b00001_000001_00001; 
		242: oled_colour = 16'b00001_000001_00001; 
		243: oled_colour = 16'b00001_000001_00001; 
		244: oled_colour = 16'b00001_000001_00001; 
		245: oled_colour = 16'b00001_000001_00001; 
		246: oled_colour = 16'b00001_000001_00001; 
		247: oled_colour = 16'b00001_000001_00001; 
		248: oled_colour = 16'b00001_000001_00001; 
		249: oled_colour = 16'b00001_000001_00001; 
		250: oled_colour = 16'b00001_000001_00001; 
		251: oled_colour = 16'b00001_000001_00001; 
		252: oled_colour = 16'b00001_000001_00001; 
		253: oled_colour = 16'b00001_000001_00001; 
		254: oled_colour = 16'b00001_000001_00001; 
		255: oled_colour = 16'b00001_000001_00001; 
		256: oled_colour = 16'b00001_000001_00001; 
		257: oled_colour = 16'b00001_000001_00001; 
		258: oled_colour = 16'b00001_000001_00001; 
		259: oled_colour = 16'b00001_000001_00001; 
		260: oled_colour = 16'b00001_000001_00001; 
		261: oled_colour = 16'b00001_000001_00001; 
		262: oled_colour = 16'b00001_000001_00001; 
		263: oled_colour = 16'b00001_000001_00001; 
		264: oled_colour = 16'b00001_000001_00001; 
		265: oled_colour = 16'b00001_000001_00001; 
		266: oled_colour = 16'b00001_000001_00001; 
		267: oled_colour = 16'b00001_000001_00001; 
		268: oled_colour = 16'b00001_000001_00001; 
		269: oled_colour = 16'b00001_000001_00001; 
		270: oled_colour = 16'b00001_000001_00001; 
		271: oled_colour = 16'b00001_000001_00001; 
		272: oled_colour = 16'b00001_000001_00001; 
		273: oled_colour = 16'b00001_000001_00001; 
		274: oled_colour = 16'b00001_000001_00001; 
		275: oled_colour = 16'b00001_000001_00001; 
		276: oled_colour = 16'b00001_000001_00001; 
		277: oled_colour = 16'b00001_000001_00001; 
		278: oled_colour = 16'b00001_000001_00001; 
		279: oled_colour = 16'b00001_000001_00001; 
		280: oled_colour = 16'b00001_000001_00001; 
		281: oled_colour = 16'b00001_000001_00001; 
		282: oled_colour = 16'b00001_000001_00001; 
		283: oled_colour = 16'b00001_000001_00001; 
		284: oled_colour = 16'b00001_000001_00001; 
		285: oled_colour = 16'b00001_000001_00001; 
		286: oled_colour = 16'b00001_000001_00001; 
		287: oled_colour = 16'b00001_000001_00001; 
		288: oled_colour = 16'b00001_000001_00001; 
		289: oled_colour = 16'b00001_000001_00001; 
		290: oled_colour = 16'b00001_000001_00001; 
		291: oled_colour = 16'b00001_000001_00001; 
		292: oled_colour = 16'b00001_000001_00001; 
		293: oled_colour = 16'b00001_000001_00001; 
		294: oled_colour = 16'b00001_000001_00001; 
		295: oled_colour = 16'b00001_000001_00001; 
		296: oled_colour = 16'b00001_000001_00001; 
		297: oled_colour = 16'b00001_000001_00001; 
		298: oled_colour = 16'b00001_000001_00001; 
		299: oled_colour = 16'b00001_000001_00001; 
		300: oled_colour = 16'b00001_000001_00001; 
		301: oled_colour = 16'b00001_000001_00001; 
		302: oled_colour = 16'b00001_000001_00001; 
		303: oled_colour = 16'b00001_000001_00001; 
		304: oled_colour = 16'b00001_000001_00001; 
		305: oled_colour = 16'b00001_000001_00001; 
		306: oled_colour = 16'b00001_000001_00001; 
		307: oled_colour = 16'b00001_000001_00001; 
		308: oled_colour = 16'b00001_000001_00001; 
		309: oled_colour = 16'b00001_000001_00001; 
		310: oled_colour = 16'b00001_000001_00001; 
		311: oled_colour = 16'b00001_000001_00001; 
		312: oled_colour = 16'b00001_000001_00001; 
		313: oled_colour = 16'b00001_000001_00001; 
		314: oled_colour = 16'b00001_000001_00001; 
		315: oled_colour = 16'b00001_000001_00001; 
		316: oled_colour = 16'b00001_000001_00001; 
		317: oled_colour = 16'b00001_000001_00001; 
		318: oled_colour = 16'b00001_000001_00001; 
		319: oled_colour = 16'b00001_000001_00001; 
		320: oled_colour = 16'b00001_000001_00001; 
		321: oled_colour = 16'b00001_000001_00001; 
		322: oled_colour = 16'b00001_000001_00001; 
		323: oled_colour = 16'b00001_000001_00001; 
		324: oled_colour = 16'b00001_000001_00001; 
		325: oled_colour = 16'b00001_000001_00001; 
		326: oled_colour = 16'b00001_000001_00001; 
		327: oled_colour = 16'b00001_000001_00001; 
		328: oled_colour = 16'b00001_000001_00001; 
		329: oled_colour = 16'b00001_000001_00001; 
		330: oled_colour = 16'b00001_000001_00001; 
		331: oled_colour = 16'b00001_000001_00001; 
		332: oled_colour = 16'b00001_000001_00001; 
		333: oled_colour = 16'b00001_000001_00001; 
		334: oled_colour = 16'b00001_000001_00001; 
		335: oled_colour = 16'b00001_000001_00001; 
		336: oled_colour = 16'b00001_000001_00001; 
		337: oled_colour = 16'b00001_000001_00001; 
		338: oled_colour = 16'b00001_000001_00001; 
		339: oled_colour = 16'b00001_000001_00001; 
		340: oled_colour = 16'b00001_000001_00001; 
		341: oled_colour = 16'b00001_000001_00001; 
		342: oled_colour = 16'b00001_000001_00001; 
		343: oled_colour = 16'b00001_000001_00001; 
		344: oled_colour = 16'b00001_000001_00001; 
		345: oled_colour = 16'b00001_000001_00001; 
		346: oled_colour = 16'b00001_000001_00001; 
		347: oled_colour = 16'b00001_000001_00001; 
		348: oled_colour = 16'b00001_000001_00001; 
		349: oled_colour = 16'b00001_000001_00001; 
		350: oled_colour = 16'b00001_000001_00001; 
		351: oled_colour = 16'b00001_000001_00001; 
		352: oled_colour = 16'b00001_000001_00001; 
		353: oled_colour = 16'b00001_000001_00001; 
		354: oled_colour = 16'b00001_000001_00001; 
		355: oled_colour = 16'b00001_000001_00001; 
		356: oled_colour = 16'b00001_000001_00001; 
		357: oled_colour = 16'b00001_000001_00001; 
		358: oled_colour = 16'b00001_000001_00001; 
		359: oled_colour = 16'b00001_000001_00001; 
		360: oled_colour = 16'b00001_000001_00001; 
		361: oled_colour = 16'b00001_000001_00001; 
		362: oled_colour = 16'b00001_000001_00001; 
		363: oled_colour = 16'b00001_000001_00001; 
		364: oled_colour = 16'b00001_000001_00001; 
		365: oled_colour = 16'b00001_000001_00001; 
		366: oled_colour = 16'b00001_000001_00001; 
		367: oled_colour = 16'b00001_000001_00001; 
		368: oled_colour = 16'b00001_000001_00001; 
		369: oled_colour = 16'b00001_000001_00001; 
		370: oled_colour = 16'b00001_000001_00001; 
		371: oled_colour = 16'b00001_000001_00001; 
		372: oled_colour = 16'b00001_000001_00001; 
		373: oled_colour = 16'b00001_000001_00001; 
		374: oled_colour = 16'b00001_000001_00001; 
		375: oled_colour = 16'b00001_000001_00001; 
		376: oled_colour = 16'b00001_000001_00001; 
		377: oled_colour = 16'b00001_000001_00001; 
		378: oled_colour = 16'b00001_000001_00001; 
		379: oled_colour = 16'b00001_000001_00001; 
		380: oled_colour = 16'b00001_000001_00001; 
		381: oled_colour = 16'b00001_000001_00001; 
		382: oled_colour = 16'b00001_000001_00001; 
		383: oled_colour = 16'b00001_000001_00001; 
		384: oled_colour = 16'b00001_000001_00001; 
		385: oled_colour = 16'b00001_000001_00001; 
		386: oled_colour = 16'b00001_000001_00001; 
		387: oled_colour = 16'b00001_000001_00001; 
		388: oled_colour = 16'b00001_000001_00001; 
		389: oled_colour = 16'b00001_000001_00001; 
		390: oled_colour = 16'b00001_000001_00001; 
		391: oled_colour = 16'b00001_000001_00001; 
		392: oled_colour = 16'b00001_000001_00001; 
		393: oled_colour = 16'b00001_000001_00001; 
		394: oled_colour = 16'b00001_000001_00001; 
		395: oled_colour = 16'b00001_000001_00001; 
		396: oled_colour = 16'b00001_000001_00001; 
		397: oled_colour = 16'b00001_000001_00001; 
		398: oled_colour = 16'b00001_000001_00001; 
		399: oled_colour = 16'b00001_000001_00001; 
		400: oled_colour = 16'b00001_000001_00001; 
		401: oled_colour = 16'b00001_000001_00001; 
		402: oled_colour = 16'b00001_000001_00001; 
		403: oled_colour = 16'b00001_000001_00001; 
		404: oled_colour = 16'b00001_000001_00001; 
		405: oled_colour = 16'b00001_000001_00001; 
		406: oled_colour = 16'b00001_000001_00001; 
		407: oled_colour = 16'b00001_000001_00001; 
		408: oled_colour = 16'b00001_000001_00001; 
		409: oled_colour = 16'b00001_000001_00001; 
		410: oled_colour = 16'b00001_000001_00001; 
		411: oled_colour = 16'b00001_000001_00001; 
		412: oled_colour = 16'b00001_000001_00001; 
		413: oled_colour = 16'b00001_000001_00001; 
		414: oled_colour = 16'b00001_000001_00001; 
		415: oled_colour = 16'b00001_000001_00001; 
		416: oled_colour = 16'b00001_000001_00001; 
		417: oled_colour = 16'b00001_000001_00001; 
		418: oled_colour = 16'b00001_000001_00001; 
		419: oled_colour = 16'b00001_000001_00001; 
		420: oled_colour = 16'b00001_000001_00001; 
		421: oled_colour = 16'b00001_000001_00001; 
		422: oled_colour = 16'b00001_000001_00001; 
		423: oled_colour = 16'b00001_000001_00001; 
		424: oled_colour = 16'b00001_000001_00001; 
		425: oled_colour = 16'b00001_000001_00001; 
		426: oled_colour = 16'b00001_000001_00001; 
		427: oled_colour = 16'b00001_000001_00001; 
		428: oled_colour = 16'b00001_000001_00001; 
		429: oled_colour = 16'b00001_000001_00001; 
		430: oled_colour = 16'b00001_000001_00001; 
		431: oled_colour = 16'b00001_000001_00001; 
		432: oled_colour = 16'b00001_000001_00001; 
		433: oled_colour = 16'b00001_000001_00001; 
		434: oled_colour = 16'b00001_000001_00001; 
		435: oled_colour = 16'b00001_000001_00001; 
		436: oled_colour = 16'b00001_000001_00001; 
		437: oled_colour = 16'b00001_000001_00001; 
		438: oled_colour = 16'b00001_000001_00001; 
		439: oled_colour = 16'b00001_000001_00001; 
		440: oled_colour = 16'b00001_000001_00001; 
		441: oled_colour = 16'b00001_000001_00001; 
		442: oled_colour = 16'b00001_000001_00001; 
		443: oled_colour = 16'b00001_000001_00001; 
		444: oled_colour = 16'b00001_000001_00001; 
		445: oled_colour = 16'b00001_000001_00001; 
		446: oled_colour = 16'b00001_000001_00001; 
		447: oled_colour = 16'b00001_000001_00001; 
		448: oled_colour = 16'b00001_000001_00001; 
		449: oled_colour = 16'b00001_000001_00001; 
		450: oled_colour = 16'b00001_000001_00001; 
		451: oled_colour = 16'b00001_000001_00001; 
		452: oled_colour = 16'b00001_000001_00001; 
		453: oled_colour = 16'b00001_000001_00001; 
		454: oled_colour = 16'b00001_000001_00001; 
		455: oled_colour = 16'b00001_000001_00001; 
		456: oled_colour = 16'b00001_000001_00001; 
		457: oled_colour = 16'b00001_000001_00001; 
		458: oled_colour = 16'b00001_000001_00001; 
		459: oled_colour = 16'b00001_000001_00001; 
		460: oled_colour = 16'b00001_000001_00001; 
		461: oled_colour = 16'b00001_000001_00001; 
		462: oled_colour = 16'b00001_000001_00001; 
		463: oled_colour = 16'b00001_000001_00001; 
		464: oled_colour = 16'b00001_000001_00001; 
		465: oled_colour = 16'b00001_000001_00001; 
		466: oled_colour = 16'b00001_000001_00001; 
		467: oled_colour = 16'b00001_000001_00001; 
		468: oled_colour = 16'b00001_000001_00001; 
		469: oled_colour = 16'b00001_000001_00001; 
		470: oled_colour = 16'b00001_000001_00001; 
		471: oled_colour = 16'b00001_000001_00001; 
		472: oled_colour = 16'b00001_000001_00001; 
		473: oled_colour = 16'b00001_000001_00001; 
		474: oled_colour = 16'b00001_000001_00001; 
		475: oled_colour = 16'b00001_000001_00001; 
		476: oled_colour = 16'b00001_000001_00001; 
		477: oled_colour = 16'b00001_000001_00001; 
		478: oled_colour = 16'b00001_000001_00001; 
		479: oled_colour = 16'b00001_000001_00001; 
		480: oled_colour = 16'b00001_000001_00001; 
		481: oled_colour = 16'b00001_000001_00001; 
		482: oled_colour = 16'b00001_000001_00001; 
		483: oled_colour = 16'b00001_000001_00001; 
		484: oled_colour = 16'b00001_000001_00001; 
		485: oled_colour = 16'b00001_000001_00001; 
		486: oled_colour = 16'b00001_000001_00001; 
		487: oled_colour = 16'b00001_000001_00001; 
		488: oled_colour = 16'b00001_000001_00001; 
		489: oled_colour = 16'b00001_000001_00001; 
		490: oled_colour = 16'b00001_000001_00001; 
		491: oled_colour = 16'b00001_000001_00001; 
		492: oled_colour = 16'b00001_000001_00001; 
		493: oled_colour = 16'b00001_000001_00001; 
		494: oled_colour = 16'b00001_000001_00001; 
		495: oled_colour = 16'b00001_000001_00001; 
		496: oled_colour = 16'b00001_000001_00001; 
		497: oled_colour = 16'b00001_000001_00001; 
		498: oled_colour = 16'b00001_000001_00001; 
		499: oled_colour = 16'b00001_000001_00001; 
		500: oled_colour = 16'b00001_000001_00001; 
		501: oled_colour = 16'b00001_000001_00001; 
		502: oled_colour = 16'b00001_000001_00001; 
		503: oled_colour = 16'b00001_000001_00001; 
		504: oled_colour = 16'b00001_000001_00001; 
		505: oled_colour = 16'b00001_000001_00001; 
		506: oled_colour = 16'b00001_000001_00001; 
		507: oled_colour = 16'b00001_000001_00001; 
		508: oled_colour = 16'b00001_000001_00001; 
		509: oled_colour = 16'b00001_000001_00001; 
		510: oled_colour = 16'b00001_000001_00001; 
		511: oled_colour = 16'b00001_000001_00001; 
		512: oled_colour = 16'b00001_000001_00001; 
		513: oled_colour = 16'b00001_000001_00001; 
		514: oled_colour = 16'b00001_000001_00001; 
		515: oled_colour = 16'b00001_000001_00001; 
		516: oled_colour = 16'b00001_000001_00001; 
		517: oled_colour = 16'b00001_000001_00001; 
		518: oled_colour = 16'b00001_000001_00001; 
		519: oled_colour = 16'b00001_000001_00001; 
		520: oled_colour = 16'b00001_000001_00001; 
		521: oled_colour = 16'b00001_000001_00001; 
		522: oled_colour = 16'b00001_000001_00001; 
		523: oled_colour = 16'b00001_000001_00001; 
		524: oled_colour = 16'b00001_000001_00001; 
		525: oled_colour = 16'b00001_000001_00001; 
		526: oled_colour = 16'b00001_000001_00001; 
		527: oled_colour = 16'b00001_000001_00001; 
		528: oled_colour = 16'b00001_000001_00001; 
		529: oled_colour = 16'b00001_000001_00001; 
		530: oled_colour = 16'b00001_000001_00001; 
		531: oled_colour = 16'b00001_000001_00001; 
		532: oled_colour = 16'b00001_000001_00001; 
		533: oled_colour = 16'b00001_000001_00001; 
		534: oled_colour = 16'b00001_000001_00001; 
		535: oled_colour = 16'b00001_000001_00001; 
		536: oled_colour = 16'b00001_000001_00001; 
		537: oled_colour = 16'b00001_000001_00001; 
		538: oled_colour = 16'b00001_000001_00001; 
		539: oled_colour = 16'b00001_000001_00001; 
		540: oled_colour = 16'b00001_000001_00001; 
		541: oled_colour = 16'b00001_000001_00001; 
		542: oled_colour = 16'b00001_000001_00001; 
		543: oled_colour = 16'b00001_000001_00001; 
		544: oled_colour = 16'b00001_000001_00001; 
		545: oled_colour = 16'b00001_000001_00001; 
		546: oled_colour = 16'b00001_000001_00001; 
		547: oled_colour = 16'b00001_000001_00001; 
		548: oled_colour = 16'b00001_000001_00001; 
		549: oled_colour = 16'b00001_000001_00001; 
		550: oled_colour = 16'b00001_000001_00001; 
		551: oled_colour = 16'b00001_000001_00001; 
		552: oled_colour = 16'b00001_000001_00001; 
		553: oled_colour = 16'b00001_000001_00001; 
		554: oled_colour = 16'b00001_000001_00001; 
		555: oled_colour = 16'b00001_000001_00001; 
		556: oled_colour = 16'b00001_000001_00001; 
		557: oled_colour = 16'b00001_000001_00001; 
		558: oled_colour = 16'b00001_000001_00001; 
		559: oled_colour = 16'b00001_000001_00001; 
		560: oled_colour = 16'b00001_000001_00001; 
		561: oled_colour = 16'b00001_000001_00001; 
		562: oled_colour = 16'b00001_000001_00001; 
		563: oled_colour = 16'b00001_000001_00001; 
		564: oled_colour = 16'b00001_000001_00001; 
		565: oled_colour = 16'b00001_000001_00001; 
		566: oled_colour = 16'b00001_000001_00001; 
		567: oled_colour = 16'b00001_000001_00001; 
		568: oled_colour = 16'b00001_000001_00001; 
		569: oled_colour = 16'b00001_000001_00001; 
		570: oled_colour = 16'b00001_000001_00001; 
		571: oled_colour = 16'b00001_000001_00001; 
		572: oled_colour = 16'b00001_000001_00001; 
		573: oled_colour = 16'b00001_000001_00001; 
		574: oled_colour = 16'b00001_000001_00001; 
		575: oled_colour = 16'b00001_000001_00001; 
		576: oled_colour = 16'b00001_000001_00001; 
		577: oled_colour = 16'b00001_000001_00001; 
		578: oled_colour = 16'b00001_000001_00001; 
		579: oled_colour = 16'b00001_000001_00001; 
		580: oled_colour = 16'b00001_000001_00001; 
		581: oled_colour = 16'b00001_000001_00001; 
		582: oled_colour = 16'b00001_000001_00001; 
		583: oled_colour = 16'b00001_000001_00001; 
		584: oled_colour = 16'b00001_000001_00001; 
		585: oled_colour = 16'b00001_000001_00001; 
		586: oled_colour = 16'b00001_000001_00001; 
		587: oled_colour = 16'b00001_000001_00001; 
		588: oled_colour = 16'b00001_000001_00001; 
		589: oled_colour = 16'b00001_000001_00001; 
		590: oled_colour = 16'b00001_000001_00001; 
		591: oled_colour = 16'b00001_000001_00001; 
		592: oled_colour = 16'b00001_000001_00001; 
		593: oled_colour = 16'b00001_000001_00001; 
		594: oled_colour = 16'b00001_000001_00001; 
		595: oled_colour = 16'b00001_000001_00001; 
		596: oled_colour = 16'b00001_000001_00001; 
		597: oled_colour = 16'b00001_000001_00001; 
		598: oled_colour = 16'b00001_000001_00001; 
		599: oled_colour = 16'b00001_000001_00001; 
		600: oled_colour = 16'b00001_000001_00001; 
		601: oled_colour = 16'b00001_000001_00001; 
		602: oled_colour = 16'b00001_000001_00001; 
		603: oled_colour = 16'b00001_000001_00001; 
		604: oled_colour = 16'b00001_000001_00001; 
		605: oled_colour = 16'b00001_000001_00001; 
		606: oled_colour = 16'b00001_000001_00001; 
		607: oled_colour = 16'b00001_000001_00001; 
		608: oled_colour = 16'b00001_000001_00001; 
		609: oled_colour = 16'b00001_000001_00001; 
		610: oled_colour = 16'b00001_000001_00001; 
		611: oled_colour = 16'b00001_000001_00001; 
		612: oled_colour = 16'b00001_000001_00001; 
		613: oled_colour = 16'b00001_000001_00001; 
		614: oled_colour = 16'b00001_000001_00001; 
		615: oled_colour = 16'b00001_000001_00001; 
		616: oled_colour = 16'b00001_000001_00001; 
		617: oled_colour = 16'b00001_000001_00001; 
		618: oled_colour = 16'b00001_000001_00001; 
		619: oled_colour = 16'b00001_000001_00001; 
		620: oled_colour = 16'b00001_000001_00001; 
		621: oled_colour = 16'b00001_000001_00001; 
		622: oled_colour = 16'b00001_000001_00001; 
		623: oled_colour = 16'b00001_000001_00001; 
		624: oled_colour = 16'b00001_000001_00001; 
		625: oled_colour = 16'b00001_000001_00001; 
		626: oled_colour = 16'b00001_000001_00001; 
		627: oled_colour = 16'b00001_000001_00001; 
		628: oled_colour = 16'b00001_000001_00001; 
		629: oled_colour = 16'b00001_000001_00001; 
		630: oled_colour = 16'b00001_000001_00001; 
		631: oled_colour = 16'b00001_000001_00001; 
		632: oled_colour = 16'b00001_000001_00001; 
		633: oled_colour = 16'b00001_000001_00001; 
		634: oled_colour = 16'b00001_000001_00001; 
		635: oled_colour = 16'b00001_000001_00001; 
		636: oled_colour = 16'b00001_000001_00001; 
		637: oled_colour = 16'b00001_000001_00001; 
		638: oled_colour = 16'b00001_000001_00001; 
		639: oled_colour = 16'b00001_000001_00001; 
		640: oled_colour = 16'b00001_000001_00001; 
		641: oled_colour = 16'b00001_000001_00001; 
		642: oled_colour = 16'b00001_000001_00001; 
		643: oled_colour = 16'b00001_000001_00001; 
		644: oled_colour = 16'b00001_000001_00001; 
		645: oled_colour = 16'b00001_000001_00001; 
		646: oled_colour = 16'b00001_000001_00001; 
		647: oled_colour = 16'b00001_000001_00001; 
		648: oled_colour = 16'b00001_000001_00001; 
		649: oled_colour = 16'b00001_000001_00001; 
		650: oled_colour = 16'b00001_000001_00001; 
		651: oled_colour = 16'b00001_000001_00001; 
		652: oled_colour = 16'b00001_000001_00001; 
		653: oled_colour = 16'b00001_000001_00001; 
		654: oled_colour = 16'b00001_000001_00001; 
		655: oled_colour = 16'b00001_000001_00001; 
		656: oled_colour = 16'b00001_000001_00001; 
		657: oled_colour = 16'b00001_000001_00001; 
		658: oled_colour = 16'b00001_000001_00001; 
		659: oled_colour = 16'b00001_000001_00001; 
		660: oled_colour = 16'b00001_000001_00001; 
		661: oled_colour = 16'b00001_000001_00001; 
		662: oled_colour = 16'b00001_000001_00001; 
		663: oled_colour = 16'b00001_000001_00001; 
		664: oled_colour = 16'b00001_000001_00001; 
		665: oled_colour = 16'b00001_000001_00001; 
		666: oled_colour = 16'b00001_000001_00001; 
		667: oled_colour = 16'b00001_000001_00001; 
		668: oled_colour = 16'b00001_000001_00001; 
		669: oled_colour = 16'b00001_000001_00001; 
		670: oled_colour = 16'b00001_000001_00001; 
		671: oled_colour = 16'b00001_000001_00001; 
		672: oled_colour = 16'b00001_000001_00001; 
		673: oled_colour = 16'b00001_000001_00001; 
		674: oled_colour = 16'b00001_000001_00001; 
		675: oled_colour = 16'b00001_000001_00001; 
		676: oled_colour = 16'b00001_000001_00001; 
		677: oled_colour = 16'b00001_000001_00001; 
		678: oled_colour = 16'b00001_000001_00001; 
		679: oled_colour = 16'b00001_000001_00001; 
		680: oled_colour = 16'b00001_000001_00001; 
		681: oled_colour = 16'b00001_000001_00001; 
		682: oled_colour = 16'b00001_000001_00001; 
		683: oled_colour = 16'b00001_000001_00001; 
		684: oled_colour = 16'b00001_000001_00001; 
		685: oled_colour = 16'b00001_000001_00001; 
		686: oled_colour = 16'b00001_000001_00001; 
		687: oled_colour = 16'b00001_000001_00001; 
		688: oled_colour = 16'b00001_000001_00001; 
		689: oled_colour = 16'b00001_000001_00001; 
		690: oled_colour = 16'b00001_000001_00001; 
		691: oled_colour = 16'b00001_000001_00001; 
		692: oled_colour = 16'b00001_000001_00001; 
		693: oled_colour = 16'b00001_000001_00001; 
		694: oled_colour = 16'b00001_000001_00001; 
		695: oled_colour = 16'b00001_000001_00001; 
		696: oled_colour = 16'b00001_000001_00001; 
		697: oled_colour = 16'b00001_000001_00001; 
		698: oled_colour = 16'b00001_000001_00001; 
		699: oled_colour = 16'b00001_000001_00001; 
		700: oled_colour = 16'b00001_000001_00001; 
		701: oled_colour = 16'b00001_000001_00001; 
		702: oled_colour = 16'b00001_000001_00001; 
		703: oled_colour = 16'b00001_000001_00001; 
		704: oled_colour = 16'b00001_000001_00001; 
		705: oled_colour = 16'b00001_000001_00001; 
		706: oled_colour = 16'b00001_000001_00001; 
		707: oled_colour = 16'b00001_000001_00001; 
		708: oled_colour = 16'b00001_000001_00001; 
		709: oled_colour = 16'b00001_000001_00001; 
		710: oled_colour = 16'b00001_000001_00001; 
		711: oled_colour = 16'b00001_000001_00001; 
		712: oled_colour = 16'b00001_000001_00001; 
		713: oled_colour = 16'b00001_000001_00001; 
		714: oled_colour = 16'b00001_000001_00001; 
		715: oled_colour = 16'b00001_000001_00001; 
		716: oled_colour = 16'b00001_000001_00001; 
		717: oled_colour = 16'b00001_000001_00001; 
		718: oled_colour = 16'b00001_000001_00001; 
		719: oled_colour = 16'b00001_000001_00001; 
		720: oled_colour = 16'b00001_000001_00001; 
		721: oled_colour = 16'b00001_000001_00001; 
		722: oled_colour = 16'b00001_000001_00001; 
		723: oled_colour = 16'b00001_000001_00001; 
		724: oled_colour = 16'b00001_000001_00001; 
		725: oled_colour = 16'b00001_000001_00001; 
		726: oled_colour = 16'b00001_000001_00001; 
		727: oled_colour = 16'b00001_000001_00001; 
		728: oled_colour = 16'b00001_000001_00001; 
		729: oled_colour = 16'b00001_000001_00001; 
		730: oled_colour = 16'b00001_000001_00001; 
		731: oled_colour = 16'b00001_000001_00001; 
		732: oled_colour = 16'b00001_000001_00001; 
		733: oled_colour = 16'b00001_000001_00001; 
		734: oled_colour = 16'b00001_000001_00001; 
		735: oled_colour = 16'b00001_000001_00001; 
		736: oled_colour = 16'b00001_000001_00001; 
		737: oled_colour = 16'b00001_000001_00001; 
		738: oled_colour = 16'b00001_000001_00001; 
		739: oled_colour = 16'b00001_000001_00001; 
		740: oled_colour = 16'b00001_000001_00001; 
		741: oled_colour = 16'b00001_000001_00001; 
		742: oled_colour = 16'b00001_000001_00001; 
		743: oled_colour = 16'b00001_000001_00001; 
		744: oled_colour = 16'b00001_000001_00001; 
		745: oled_colour = 16'b00001_000001_00001; 
		746: oled_colour = 16'b00001_000001_00001; 
		747: oled_colour = 16'b00001_000001_00001; 
		748: oled_colour = 16'b00001_000001_00001; 
		749: oled_colour = 16'b00001_000001_00001; 
		750: oled_colour = 16'b00001_000001_00001; 
		751: oled_colour = 16'b00001_000001_00001; 
		752: oled_colour = 16'b00001_000001_00001; 
		753: oled_colour = 16'b00001_000001_00001; 
		754: oled_colour = 16'b00001_000001_00001; 
		755: oled_colour = 16'b00001_000001_00001; 
		756: oled_colour = 16'b00001_000001_00001; 
		757: oled_colour = 16'b00001_000001_00001; 
		758: oled_colour = 16'b00001_000001_00001; 
		759: oled_colour = 16'b00001_000001_00001; 
		760: oled_colour = 16'b00001_000001_00001; 
		761: oled_colour = 16'b00001_000001_00001; 
		762: oled_colour = 16'b00001_000001_00001; 
		763: oled_colour = 16'b00001_000001_00001; 
		764: oled_colour = 16'b00001_000001_00001; 
		765: oled_colour = 16'b00001_000001_00001; 
		766: oled_colour = 16'b00001_000001_00001; 
		767: oled_colour = 16'b00001_000001_00001; 
		768: oled_colour = 16'b00001_000001_00001; 
		769: oled_colour = 16'b00001_000001_00001; 
		770: oled_colour = 16'b00001_000001_00001; 
		771: oled_colour = 16'b00001_000001_00001; 
		772: oled_colour = 16'b00001_000001_00001; 
		773: oled_colour = 16'b00001_000001_00001; 
		774: oled_colour = 16'b00001_000001_00001; 
		775: oled_colour = 16'b00001_000001_00001; 
		776: oled_colour = 16'b00001_000001_00001; 
		777: oled_colour = 16'b00001_000001_00001; 
		778: oled_colour = 16'b00001_000001_00001; 
		779: oled_colour = 16'b00001_000001_00001; 
		780: oled_colour = 16'b00001_000001_00001; 
		781: oled_colour = 16'b00001_000001_00001; 
		782: oled_colour = 16'b00001_000001_00001; 
		783: oled_colour = 16'b00001_000001_00001; 
		784: oled_colour = 16'b00001_000001_00001; 
		785: oled_colour = 16'b00001_000001_00001; 
		786: oled_colour = 16'b00001_000001_00001; 
		787: oled_colour = 16'b00001_000001_00001; 
		788: oled_colour = 16'b00001_000001_00001; 
		789: oled_colour = 16'b00001_000001_00001; 
		790: oled_colour = 16'b00001_000001_00001; 
		791: oled_colour = 16'b00001_000001_00001; 
		792: oled_colour = 16'b00001_000001_00001; 
		793: oled_colour = 16'b00001_000001_00001; 
		794: oled_colour = 16'b00001_000001_00001; 
		795: oled_colour = 16'b00001_000001_00001; 
		796: oled_colour = 16'b00001_000001_00001; 
		797: oled_colour = 16'b00001_000001_00001; 
		798: oled_colour = 16'b00001_000001_00001; 
		799: oled_colour = 16'b00001_000001_00001; 
		800: oled_colour = 16'b00001_000001_00001; 
		801: oled_colour = 16'b00001_000001_00001; 
		802: oled_colour = 16'b00001_000001_00001; 
		803: oled_colour = 16'b00001_000001_00001; 
		804: oled_colour = 16'b00001_000001_00001; 
		805: oled_colour = 16'b00001_000001_00001; 
		806: oled_colour = 16'b00001_000001_00001; 
		807: oled_colour = 16'b00001_000001_00001; 
		808: oled_colour = 16'b00001_000001_00001; 
		809: oled_colour = 16'b00001_000001_00001; 
		810: oled_colour = 16'b00001_000001_00001; 
		811: oled_colour = 16'b00001_000001_00001; 
		812: oled_colour = 16'b00001_000001_00001; 
		813: oled_colour = 16'b00001_000001_00001; 
		814: oled_colour = 16'b00001_000001_00001; 
		815: oled_colour = 16'b00001_000001_00001; 
		816: oled_colour = 16'b00001_000001_00001; 
		817: oled_colour = 16'b00001_000001_00001; 
		818: oled_colour = 16'b00001_000001_00001; 
		819: oled_colour = 16'b00001_000001_00001; 
		820: oled_colour = 16'b00001_000001_00001; 
		821: oled_colour = 16'b00001_000001_00001; 
		822: oled_colour = 16'b00001_000001_00001; 
		823: oled_colour = 16'b00001_000001_00001; 
		824: oled_colour = 16'b00001_000001_00001; 
		825: oled_colour = 16'b00001_000001_00001; 
		826: oled_colour = 16'b00001_000001_00001; 
		827: oled_colour = 16'b00001_000001_00001; 
		828: oled_colour = 16'b00001_000001_00001; 
		829: oled_colour = 16'b00001_000001_00001; 
		830: oled_colour = 16'b00001_000001_00001; 
		831: oled_colour = 16'b00001_000001_00001; 
		832: oled_colour = 16'b00001_000001_00001; 
		833: oled_colour = 16'b00001_000001_00001; 
		834: oled_colour = 16'b00001_000001_00001; 
		835: oled_colour = 16'b00001_000001_00001; 
		836: oled_colour = 16'b00001_000001_00001; 
		837: oled_colour = 16'b00001_000001_00001; 
		838: oled_colour = 16'b00001_000001_00001; 
		839: oled_colour = 16'b00001_000001_00001; 
		840: oled_colour = 16'b00001_000001_00001; 
		841: oled_colour = 16'b00001_000001_00001; 
		842: oled_colour = 16'b00001_000001_00001; 
		843: oled_colour = 16'b00001_000001_00001; 
		844: oled_colour = 16'b00001_000001_00001; 
		845: oled_colour = 16'b00001_000001_00001; 
		846: oled_colour = 16'b00001_000001_00001; 
		847: oled_colour = 16'b00001_000001_00001; 
		848: oled_colour = 16'b00001_000001_00001; 
		849: oled_colour = 16'b00001_000001_00001; 
		850: oled_colour = 16'b00001_000001_00001; 
		851: oled_colour = 16'b00001_000001_00001; 
		852: oled_colour = 16'b00001_000001_00001; 
		853: oled_colour = 16'b00001_000001_00001; 
		854: oled_colour = 16'b00001_000001_00001; 
		855: oled_colour = 16'b00001_000001_00001; 
		856: oled_colour = 16'b00001_000001_00001; 
		857: oled_colour = 16'b00001_000001_00001; 
		858: oled_colour = 16'b00001_000001_00001; 
		859: oled_colour = 16'b00001_000001_00001; 
		860: oled_colour = 16'b00001_000001_00001; 
		861: oled_colour = 16'b00001_000001_00001; 
		862: oled_colour = 16'b00001_000001_00001; 
		863: oled_colour = 16'b00001_000001_00001; 
		864: oled_colour = 16'b00001_000001_00001; 
		865: oled_colour = 16'b00001_000001_00001; 
		866: oled_colour = 16'b00001_000001_00001; 
		867: oled_colour = 16'b00001_000001_00001; 
		868: oled_colour = 16'b00001_000001_00001; 
		869: oled_colour = 16'b00001_000001_00001; 
		870: oled_colour = 16'b00001_000001_00001; 
		871: oled_colour = 16'b00001_000001_00001; 
		872: oled_colour = 16'b00001_000001_00001; 
		873: oled_colour = 16'b00001_000001_00001; 
		874: oled_colour = 16'b00001_000001_00001; 
		875: oled_colour = 16'b00001_000001_00001; 
		876: oled_colour = 16'b00001_000001_00001; 
		877: oled_colour = 16'b00001_000001_00001; 
		878: oled_colour = 16'b00001_000001_00001; 
		879: oled_colour = 16'b00001_000001_00001; 
		880: oled_colour = 16'b00001_000001_00001; 
		881: oled_colour = 16'b00001_000001_00001; 
		882: oled_colour = 16'b00001_000001_00001; 
		883: oled_colour = 16'b00001_000001_00001; 
		884: oled_colour = 16'b00001_000001_00001; 
		885: oled_colour = 16'b00001_000001_00001; 
		886: oled_colour = 16'b00001_000001_00001; 
		887: oled_colour = 16'b00001_000001_00001; 
		888: oled_colour = 16'b00001_000001_00001; 
		889: oled_colour = 16'b00001_000001_00001; 
		890: oled_colour = 16'b00001_000001_00001; 
		891: oled_colour = 16'b00001_000001_00001; 
		892: oled_colour = 16'b00001_000001_00001; 
		893: oled_colour = 16'b00001_000001_00001; 
		894: oled_colour = 16'b00001_000001_00001; 
		895: oled_colour = 16'b00001_000001_00001; 
		896: oled_colour = 16'b00001_000001_00001; 
		897: oled_colour = 16'b00001_000001_00001; 
		898: oled_colour = 16'b00001_000001_00001; 
		899: oled_colour = 16'b00001_000001_00001; 
		900: oled_colour = 16'b00001_000001_00001; 
		901: oled_colour = 16'b00001_000001_00001; 
		902: oled_colour = 16'b00001_000001_00001; 
		903: oled_colour = 16'b00001_000001_00001; 
		904: oled_colour = 16'b00001_000001_00001; 
		905: oled_colour = 16'b00001_000001_00001; 
		906: oled_colour = 16'b00001_000001_00001; 
		907: oled_colour = 16'b00001_000001_00001; 
		908: oled_colour = 16'b00001_000001_00001; 
		909: oled_colour = 16'b00001_000001_00001; 
		910: oled_colour = 16'b00001_000001_00001; 
		911: oled_colour = 16'b00001_000001_00001; 
		912: oled_colour = 16'b00001_000001_00001; 
		913: oled_colour = 16'b00001_000001_00001; 
		914: oled_colour = 16'b00001_000001_00001; 
		915: oled_colour = 16'b00001_000001_00001; 
		916: oled_colour = 16'b00001_000001_00001; 
		917: oled_colour = 16'b00001_000001_00001; 
		918: oled_colour = 16'b00001_000001_00001; 
		919: oled_colour = 16'b00001_000001_00001; 
		920: oled_colour = 16'b00001_000001_00001; 
		921: oled_colour = 16'b00001_000001_00001; 
		922: oled_colour = 16'b00001_000001_00001; 
		923: oled_colour = 16'b00001_000001_00001; 
		924: oled_colour = 16'b00001_000001_00001; 
		925: oled_colour = 16'b00001_000001_00001; 
		926: oled_colour = 16'b00001_000001_00001; 
		927: oled_colour = 16'b00001_000001_00001; 
		928: oled_colour = 16'b00001_000001_00001; 
		929: oled_colour = 16'b00001_000001_00001; 
		930: oled_colour = 16'b00001_000001_00001; 
		931: oled_colour = 16'b00001_000001_00001; 
		932: oled_colour = 16'b00001_000001_00001; 
		933: oled_colour = 16'b00001_000001_00001; 
		934: oled_colour = 16'b00001_000001_00001; 
		935: oled_colour = 16'b00001_000001_00001; 
		936: oled_colour = 16'b00001_000001_00001; 
		937: oled_colour = 16'b00001_000001_00001; 
		938: oled_colour = 16'b00001_000001_00001; 
		939: oled_colour = 16'b00001_000001_00001; 
		940: oled_colour = 16'b00001_000001_00001; 
		941: oled_colour = 16'b00001_000001_00001; 
		942: oled_colour = 16'b00001_000001_00001; 
		943: oled_colour = 16'b00001_000001_00001; 
		944: oled_colour = 16'b00001_000001_00001; 
		945: oled_colour = 16'b00001_000001_00001; 
		946: oled_colour = 16'b00001_000001_00001; 
		947: oled_colour = 16'b00001_000001_00001; 
		948: oled_colour = 16'b00001_000001_00001; 
		949: oled_colour = 16'b00001_000001_00001; 
		950: oled_colour = 16'b00001_000001_00001; 
		951: oled_colour = 16'b00001_000001_00001; 
		952: oled_colour = 16'b00001_000001_00001; 
		953: oled_colour = 16'b00001_000001_00001; 
		954: oled_colour = 16'b00001_000001_00001; 
		955: oled_colour = 16'b00001_000001_00001; 
		956: oled_colour = 16'b00001_000001_00001; 
		957: oled_colour = 16'b00001_000001_00001; 
		958: oled_colour = 16'b00001_000001_00001; 
		959: oled_colour = 16'b00001_000001_00001; 
		960: oled_colour = 16'b00001_000001_00001; 
		961: oled_colour = 16'b00001_000001_00001; 
		962: oled_colour = 16'b00001_000001_00001; 
		963: oled_colour = 16'b00001_000001_00001; 
		964: oled_colour = 16'b00001_000001_00001; 
		965: oled_colour = 16'b00001_000001_00001; 
		966: oled_colour = 16'b00001_000001_00001; 
		967: oled_colour = 16'b00001_000001_00001; 
		968: oled_colour = 16'b00001_000001_00001; 
		969: oled_colour = 16'b00001_000001_00001; 
		970: oled_colour = 16'b00001_000001_00001; 
		971: oled_colour = 16'b00001_000001_00001; 
		972: oled_colour = 16'b00001_000001_00001; 
		973: oled_colour = 16'b00001_000001_00001; 
		974: oled_colour = 16'b00001_000001_00001; 
		975: oled_colour = 16'b00001_000001_00001; 
		976: oled_colour = 16'b00001_000001_00001; 
		977: oled_colour = 16'b00001_000001_00001; 
		978: oled_colour = 16'b00001_000001_00001; 
		979: oled_colour = 16'b00001_000001_00001; 
		980: oled_colour = 16'b00001_000001_00001; 
		981: oled_colour = 16'b00001_000001_00001; 
		982: oled_colour = 16'b00001_000001_00001; 
		983: oled_colour = 16'b00001_000001_00001; 
		984: oled_colour = 16'b00001_000001_00001; 
		985: oled_colour = 16'b00001_000001_00001; 
		986: oled_colour = 16'b00001_000001_00001; 
		987: oled_colour = 16'b00001_000001_00001; 
		988: oled_colour = 16'b00001_000001_00001; 
		989: oled_colour = 16'b00001_000001_00001; 
		990: oled_colour = 16'b00001_000001_00001; 
		991: oled_colour = 16'b00001_000001_00001; 
		992: oled_colour = 16'b00001_000001_00001; 
		993: oled_colour = 16'b00001_000001_00001; 
		994: oled_colour = 16'b00001_000001_00001; 
		995: oled_colour = 16'b00001_000001_00001; 
		996: oled_colour = 16'b00001_000001_00001; 
		997: oled_colour = 16'b00001_000001_00001; 
		998: oled_colour = 16'b00001_000001_00001; 
		999: oled_colour = 16'b00001_000001_00001; 
		1000: oled_colour = 16'b00001_000001_00001; 
		1001: oled_colour = 16'b00001_000001_00001; 
		1002: oled_colour = 16'b00001_000001_00001; 
		1003: oled_colour = 16'b00001_000001_00001; 
		1004: oled_colour = 16'b00001_000001_00001; 
		1005: oled_colour = 16'b00001_000001_00001; 
		1006: oled_colour = 16'b00001_000001_00001; 
		1007: oled_colour = 16'b00001_000001_00001; 
		1008: oled_colour = 16'b00001_000001_00001; 
		1009: oled_colour = 16'b00001_000001_00001; 
		1010: oled_colour = 16'b00001_000001_00001; 
		1011: oled_colour = 16'b00001_000001_00001; 
		1012: oled_colour = 16'b00001_000001_00001; 
		1013: oled_colour = 16'b00001_000001_00001; 
		1014: oled_colour = 16'b00001_000001_00001; 
		1015: oled_colour = 16'b00001_000001_00001; 
		1016: oled_colour = 16'b00001_000001_00001; 
		1017: oled_colour = 16'b00001_000001_00001; 
		1018: oled_colour = 16'b00001_000001_00001; 
		1019: oled_colour = 16'b00001_000001_00001; 
		1020: oled_colour = 16'b00001_000001_00001; 
		1021: oled_colour = 16'b00001_000001_00001; 
		1022: oled_colour = 16'b00001_000001_00001; 
		1023: oled_colour = 16'b00001_000001_00001; 
		1024: oled_colour = 16'b00001_000001_00001; 
		1025: oled_colour = 16'b00001_000001_00001; 
		1026: oled_colour = 16'b00001_000001_00001; 
		1027: oled_colour = 16'b00001_000001_00001; 
		1028: oled_colour = 16'b00001_000001_00001; 
		1029: oled_colour = 16'b00001_000001_00001; 
		1030: oled_colour = 16'b00001_000001_00001; 
		1031: oled_colour = 16'b00001_000001_00001; 
		1032: oled_colour = 16'b00001_000001_00001; 
		1033: oled_colour = 16'b00001_000001_00001; 
		1034: oled_colour = 16'b00001_000001_00001; 
		1035: oled_colour = 16'b00001_000001_00001; 
		1036: oled_colour = 16'b00001_000001_00001; 
		1037: oled_colour = 16'b00001_000001_00001; 
		1038: oled_colour = 16'b00001_000001_00001; 
		1039: oled_colour = 16'b00001_000001_00001; 
		1040: oled_colour = 16'b00001_000001_00001; 
		1041: oled_colour = 16'b00001_000001_00001; 
		1042: oled_colour = 16'b00001_000001_00001; 
		1043: oled_colour = 16'b00001_000001_00001; 
		1044: oled_colour = 16'b00001_000001_00001; 
		1045: oled_colour = 16'b00001_000001_00001; 
		1046: oled_colour = 16'b00001_000001_00001; 
		1047: oled_colour = 16'b00001_000001_00001; 
		1048: oled_colour = 16'b00001_000001_00001; 
		1049: oled_colour = 16'b00001_000001_00001; 
		1050: oled_colour = 16'b00001_000001_00001; 
		1051: oled_colour = 16'b00001_000001_00001; 
		1052: oled_colour = 16'b00001_000001_00001; 
		1053: oled_colour = 16'b00001_000001_00001; 
		1054: oled_colour = 16'b00001_000001_00001; 
		1055: oled_colour = 16'b00001_000001_00001; 
		1056: oled_colour = 16'b00001_000001_00001; 
		1057: oled_colour = 16'b00001_000001_00001; 
		1058: oled_colour = 16'b00001_000001_00001; 
		1059: oled_colour = 16'b00001_000001_00001; 
		1060: oled_colour = 16'b00001_000001_00001; 
		1061: oled_colour = 16'b00001_000001_00001; 
		1062: oled_colour = 16'b00001_000001_00001; 
		1063: oled_colour = 16'b00001_000001_00001; 
		1064: oled_colour = 16'b00001_000001_00001; 
		1065: oled_colour = 16'b00001_000001_00001; 
		1066: oled_colour = 16'b00001_000001_00001; 
		1067: oled_colour = 16'b00001_000001_00001; 
		1068: oled_colour = 16'b00001_000001_00001; 
		1069: oled_colour = 16'b00001_000001_00001; 
		1070: oled_colour = 16'b00001_000001_00001; 
		1071: oled_colour = 16'b00001_000001_00001; 
		1072: oled_colour = 16'b00001_000001_00001; 
		1073: oled_colour = 16'b00001_000001_00001; 
		1074: oled_colour = 16'b00001_000001_00001; 
		1075: oled_colour = 16'b00001_000001_00001; 
		1076: oled_colour = 16'b00001_000001_00001; 
		1077: oled_colour = 16'b00001_000001_00001; 
		1078: oled_colour = 16'b00001_000001_00001; 
		1079: oled_colour = 16'b00001_000001_00001; 
		1080: oled_colour = 16'b00001_000001_00001; 
		1081: oled_colour = 16'b00001_000001_00001; 
		1082: oled_colour = 16'b00001_000001_00001; 
		1083: oled_colour = 16'b00001_000001_00001; 
		1084: oled_colour = 16'b00001_000001_00001; 
		1085: oled_colour = 16'b00001_000001_00001; 
		1086: oled_colour = 16'b00001_000001_00001; 
		1087: oled_colour = 16'b00001_000001_00001; 
		1088: oled_colour = 16'b00001_000001_00001; 
		1089: oled_colour = 16'b00001_000001_00001; 
		1090: oled_colour = 16'b00001_000001_00001; 
		1091: oled_colour = 16'b00001_000001_00001; 
		1092: oled_colour = 16'b00001_000001_00001; 
		1093: oled_colour = 16'b00001_000001_00001; 
		1094: oled_colour = 16'b00001_000001_00001; 
		1095: oled_colour = 16'b00001_000001_00001; 
		1096: oled_colour = 16'b00001_000001_00001; 
		1097: oled_colour = 16'b00001_000001_00001; 
		1098: oled_colour = 16'b00001_000001_00001; 
		1099: oled_colour = 16'b00001_000001_00001; 
		1100: oled_colour = 16'b00001_000001_00001; 
		1101: oled_colour = 16'b00001_000001_00001; 
		1102: oled_colour = 16'b00001_000001_00001; 
		1103: oled_colour = 16'b00001_000001_00001; 
		1104: oled_colour = 16'b00001_000001_00001; 
		1105: oled_colour = 16'b00001_000001_00001; 
		1106: oled_colour = 16'b00001_000001_00001; 
		1107: oled_colour = 16'b00001_000001_00001; 
		1108: oled_colour = 16'b00001_000001_00001; 
		1109: oled_colour = 16'b00001_000001_00001; 
		1110: oled_colour = 16'b00001_000001_00001; 
		1111: oled_colour = 16'b00001_000001_00001; 
		1112: oled_colour = 16'b00001_000001_00001; 
		1113: oled_colour = 16'b00001_000001_00001; 
		1114: oled_colour = 16'b00001_000001_00001; 
		1115: oled_colour = 16'b00001_000001_00001; 
		1116: oled_colour = 16'b00001_000001_00001; 
		1117: oled_colour = 16'b00001_000001_00001; 
		1118: oled_colour = 16'b00001_000001_00001; 
		1119: oled_colour = 16'b00001_000001_00001; 
		1120: oled_colour = 16'b00001_000001_00001; 
		1121: oled_colour = 16'b00001_000001_00001; 
		1122: oled_colour = 16'b00001_000001_00001; 
		1123: oled_colour = 16'b00001_000001_00001; 
		1124: oled_colour = 16'b00001_000001_00001; 
		1125: oled_colour = 16'b00001_000001_00001; 
		1126: oled_colour = 16'b00001_000001_00001; 
		1127: oled_colour = 16'b00001_000001_00001; 
		1128: oled_colour = 16'b00001_000001_00001; 
		1129: oled_colour = 16'b00001_000001_00001; 
		1130: oled_colour = 16'b00001_000001_00001; 
		1131: oled_colour = 16'b00001_000001_00001; 
		1132: oled_colour = 16'b00001_000001_00001; 
		1133: oled_colour = 16'b00001_000001_00001; 
		1134: oled_colour = 16'b00001_000001_00001; 
		1135: oled_colour = 16'b00001_000001_00001; 
		1136: oled_colour = 16'b00001_000001_00001; 
		1137: oled_colour = 16'b00001_000001_00001; 
		1138: oled_colour = 16'b00001_000001_00001; 
		1139: oled_colour = 16'b00001_000001_00001; 
		1140: oled_colour = 16'b00001_000001_00001; 
		1141: oled_colour = 16'b00001_000001_00001; 
		1142: oled_colour = 16'b00001_000001_00001; 
		1143: oled_colour = 16'b00001_000001_00001; 
		1144: oled_colour = 16'b00001_000001_00001; 
		1145: oled_colour = 16'b00001_000001_00001; 
		1146: oled_colour = 16'b00001_000001_00001; 
		1147: oled_colour = 16'b00001_000001_00001; 
		1148: oled_colour = 16'b00001_000001_00001; 
		1149: oled_colour = 16'b00001_000001_00001; 
		1150: oled_colour = 16'b00001_000001_00001; 
		1151: oled_colour = 16'b00001_000001_00001; 
		1152: oled_colour = 16'b00001_000001_00001; 
		1153: oled_colour = 16'b00001_000001_00001; 
		1154: oled_colour = 16'b00001_000001_00001; 
		1155: oled_colour = 16'b00001_000001_00001; 
		1156: oled_colour = 16'b00001_000001_00001; 
		1157: oled_colour = 16'b00001_000001_00001; 
		1158: oled_colour = 16'b00001_000001_00001; 
		1159: oled_colour = 16'b00001_000001_00001; 
		1160: oled_colour = 16'b00001_000001_00001; 
		1161: oled_colour = 16'b00001_000001_00001; 
		1162: oled_colour = 16'b00001_000001_00001; 
		1163: oled_colour = 16'b00001_000001_00001; 
		1164: oled_colour = 16'b00001_000001_00001; 
		1165: oled_colour = 16'b00001_000001_00001; 
		1166: oled_colour = 16'b00001_000001_00001; 
		1167: oled_colour = 16'b00001_000001_00001; 
		1168: oled_colour = 16'b00001_000001_00001; 
		1169: oled_colour = 16'b00001_000001_00001; 
		1170: oled_colour = 16'b00001_000001_00001; 
		1171: oled_colour = 16'b00001_000001_00001; 
		1172: oled_colour = 16'b00001_000001_00001; 
		1173: oled_colour = 16'b00001_000001_00001; 
		1174: oled_colour = 16'b00001_000001_00001; 
		1175: oled_colour = 16'b00001_000001_00001; 
		1176: oled_colour = 16'b00001_000001_00001; 
		1177: oled_colour = 16'b00001_000001_00001; 
		1178: oled_colour = 16'b00001_000001_00001; 
		1179: oled_colour = 16'b00001_000001_00001; 
		1180: oled_colour = 16'b00001_000001_00001; 
		1181: oled_colour = 16'b00001_000001_00001; 
		1182: oled_colour = 16'b00001_000001_00001; 
		1183: oled_colour = 16'b00001_000001_00001; 
		1184: oled_colour = 16'b00001_000001_00001; 
		1185: oled_colour = 16'b00001_000001_00001; 
		1186: oled_colour = 16'b00001_000001_00001; 
		1187: oled_colour = 16'b00001_000001_00001; 
		1188: oled_colour = 16'b00001_000001_00001; 
		1189: oled_colour = 16'b00001_000001_00001; 
		1190: oled_colour = 16'b00001_000001_00001; 
		1191: oled_colour = 16'b00001_000001_00001; 
		1192: oled_colour = 16'b00001_000001_00001; 
		1193: oled_colour = 16'b00001_000001_00001; 
		1194: oled_colour = 16'b00001_000001_00001; 
		1195: oled_colour = 16'b00001_000001_00001; 
		1196: oled_colour = 16'b00001_000001_00001; 
		1197: oled_colour = 16'b00001_000001_00001; 
		1198: oled_colour = 16'b00001_000001_00001; 
		1199: oled_colour = 16'b00001_000001_00001; 
		1200: oled_colour = 16'b00001_000001_00001; 
		1201: oled_colour = 16'b00001_000001_00001; 
		1202: oled_colour = 16'b00001_000001_00001; 
		1203: oled_colour = 16'b00001_000001_00001; 
		1204: oled_colour = 16'b00001_000001_00001; 
		1205: oled_colour = 16'b00001_000001_00001; 
		1206: oled_colour = 16'b00001_000001_00001; 
		1207: oled_colour = 16'b00001_000001_00001; 
		1208: oled_colour = 16'b00001_000001_00001; 
		1209: oled_colour = 16'b00001_000001_00001; 
		1210: oled_colour = 16'b00001_000001_00001; 
		1211: oled_colour = 16'b00001_000001_00001; 
		1212: oled_colour = 16'b00001_000001_00001; 
		1213: oled_colour = 16'b00001_000001_00001; 
		1214: oled_colour = 16'b00001_000001_00001; 
		1215: oled_colour = 16'b00001_000001_00001; 
		1216: oled_colour = 16'b00001_000001_00001; 
		1217: oled_colour = 16'b00001_000001_00001; 
		1218: oled_colour = 16'b00001_000001_00001; 
		1219: oled_colour = 16'b00001_000001_00001; 
		1220: oled_colour = 16'b00001_000001_00001; 
		1221: oled_colour = 16'b00001_000001_00001; 
		1222: oled_colour = 16'b00001_000001_00001; 
		1223: oled_colour = 16'b00001_000001_00001; 
		1224: oled_colour = 16'b00001_000001_00001; 
		1225: oled_colour = 16'b00001_000001_00001; 
		1226: oled_colour = 16'b00001_000001_00001; 
		1227: oled_colour = 16'b00001_000001_00001; 
		1228: oled_colour = 16'b00001_000001_00001; 
		1229: oled_colour = 16'b00001_000001_00001; 
		1230: oled_colour = 16'b00001_000001_00001; 
		1231: oled_colour = 16'b00001_000001_00001; 
		1232: oled_colour = 16'b00001_000001_00001; 
		1233: oled_colour = 16'b00001_000001_00001; 
		1234: oled_colour = 16'b00001_000001_00001; 
		1235: oled_colour = 16'b00001_000001_00001; 
		1236: oled_colour = 16'b00001_000001_00001; 
		1237: oled_colour = 16'b00001_000001_00001; 
		1238: oled_colour = 16'b00001_000001_00001; 
		1239: oled_colour = 16'b00001_000001_00001; 
		1240: oled_colour = 16'b00001_000001_00001; 
		1241: oled_colour = 16'b00001_000001_00001; 
		1242: oled_colour = 16'b00001_000001_00001; 
		1243: oled_colour = 16'b00001_000001_00001; 
		1244: oled_colour = 16'b00001_000001_00001; 
		1245: oled_colour = 16'b00001_000001_00001; 
		1246: oled_colour = 16'b00001_000001_00001; 
		1247: oled_colour = 16'b00001_000001_00001; 
		1248: oled_colour = 16'b00001_000001_00001; 
		1249: oled_colour = 16'b00001_000001_00001; 
		1250: oled_colour = 16'b00001_000001_00001; 
		1251: oled_colour = 16'b00001_000001_00001; 
		1252: oled_colour = 16'b00001_000001_00001; 
		1253: oled_colour = 16'b00001_000001_00001; 
		1254: oled_colour = 16'b00001_000001_00001; 
		1255: oled_colour = 16'b00001_000001_00001; 
		1256: oled_colour = 16'b00001_000001_00001; 
		1257: oled_colour = 16'b00001_000001_00001; 
		1258: oled_colour = 16'b00001_000001_00001; 
		1259: oled_colour = 16'b00001_000001_00001; 
		1260: oled_colour = 16'b00001_000001_00001; 
		1261: oled_colour = 16'b00001_000001_00001; 
		1262: oled_colour = 16'b00001_000001_00001; 
		1263: oled_colour = 16'b00001_000001_00001; 
		1264: oled_colour = 16'b00001_000001_00001; 
		1265: oled_colour = 16'b00001_000001_00001; 
		1266: oled_colour = 16'b00001_000001_00001; 
		1267: oled_colour = 16'b00001_000001_00001; 
		1268: oled_colour = 16'b00001_000001_00001; 
		1269: oled_colour = 16'b00001_000001_00001; 
		1270: oled_colour = 16'b00001_000001_00001; 
		1271: oled_colour = 16'b00001_000001_00001; 
		1272: oled_colour = 16'b00001_000001_00001; 
		1273: oled_colour = 16'b00001_000001_00001; 
		1274: oled_colour = 16'b00001_000001_00001; 
		1275: oled_colour = 16'b00001_000001_00001; 
		1276: oled_colour = 16'b00001_000001_00001; 
		1277: oled_colour = 16'b00001_000001_00001; 
		1278: oled_colour = 16'b00001_000001_00001; 
		1279: oled_colour = 16'b00001_000001_00001; 
		1280: oled_colour = 16'b00001_000001_00001; 
		1281: oled_colour = 16'b00001_000001_00001; 
		1282: oled_colour = 16'b00001_000001_00001; 
		1283: oled_colour = 16'b00001_000001_00001; 
		1284: oled_colour = 16'b00001_000001_00001; 
		1285: oled_colour = 16'b00001_000001_00001; 
		1286: oled_colour = 16'b00001_000001_00001; 
		1287: oled_colour = 16'b00001_000001_00001; 
		1288: oled_colour = 16'b00001_000001_00001; 
		1289: oled_colour = 16'b00001_000001_00001; 
		1290: oled_colour = 16'b00001_000001_00001; 
		1291: oled_colour = 16'b00001_000001_00001; 
		1292: oled_colour = 16'b00001_000001_00001; 
		1293: oled_colour = 16'b00001_000001_00001; 
		1294: oled_colour = 16'b00001_000001_00001; 
		1295: oled_colour = 16'b00001_000001_00001; 
		1296: oled_colour = 16'b00001_000001_00001; 
		1297: oled_colour = 16'b00001_000001_00001; 
		1298: oled_colour = 16'b00001_000001_00001; 
		1299: oled_colour = 16'b00001_000001_00001; 
		1300: oled_colour = 16'b00001_000001_00001; 
		1301: oled_colour = 16'b00001_000001_00001; 
		1302: oled_colour = 16'b00001_000001_00001; 
		1303: oled_colour = 16'b00001_000001_00001; 
		1304: oled_colour = 16'b00001_000001_00001; 
		1305: oled_colour = 16'b00001_000001_00001; 
		1306: oled_colour = 16'b00001_000001_00001; 
		1307: oled_colour = 16'b00001_000001_00001; 
		1308: oled_colour = 16'b00001_000001_00001; 
		1309: oled_colour = 16'b00001_000001_00001; 
		1310: oled_colour = 16'b00001_000001_00001; 
		1311: oled_colour = 16'b00001_000001_00001; 
		1312: oled_colour = 16'b00001_000001_00001; 
		1313: oled_colour = 16'b00001_000001_00001; 
		1314: oled_colour = 16'b00001_000001_00001; 
		1315: oled_colour = 16'b00001_000001_00001; 
		1316: oled_colour = 16'b00001_000001_00001; 
		1317: oled_colour = 16'b00001_000001_00001; 
		1318: oled_colour = 16'b00001_000001_00001; 
		1319: oled_colour = 16'b00001_000001_00001; 
		1320: oled_colour = 16'b00001_000001_00001; 
		1321: oled_colour = 16'b00001_000001_00001; 
		1322: oled_colour = 16'b00001_000001_00001; 
		1323: oled_colour = 16'b00001_000001_00001; 
		1324: oled_colour = 16'b00001_000001_00001; 
		1325: oled_colour = 16'b00001_000001_00001; 
		1326: oled_colour = 16'b00001_000001_00001; 
		1327: oled_colour = 16'b00001_000001_00001; 
		1328: oled_colour = 16'b00001_000001_00001; 
		1329: oled_colour = 16'b00001_000001_00001; 
		1330: oled_colour = 16'b00001_000001_00001; 
		1331: oled_colour = 16'b00001_000001_00001; 
		1332: oled_colour = 16'b00001_000001_00001; 
		1333: oled_colour = 16'b00001_000001_00001; 
		1334: oled_colour = 16'b00001_000001_00001; 
		1335: oled_colour = 16'b00001_000001_00001; 
		1336: oled_colour = 16'b00001_000001_00001; 
		1337: oled_colour = 16'b00001_000001_00001; 
		1338: oled_colour = 16'b00001_000001_00001; 
		1339: oled_colour = 16'b00001_000001_00001; 
		1340: oled_colour = 16'b00001_000001_00001; 
		1341: oled_colour = 16'b00001_000001_00001; 
		1342: oled_colour = 16'b00001_000001_00001; 
		1343: oled_colour = 16'b00001_000001_00001; 
		1344: oled_colour = 16'b00001_000001_00001; 
		1345: oled_colour = 16'b00001_000001_00001; 
		1346: oled_colour = 16'b00001_000001_00001; 
		1347: oled_colour = 16'b00001_000001_00001; 
		1348: oled_colour = 16'b00001_000001_00001; 
		1349: oled_colour = 16'b00001_000001_00001; 
		1350: oled_colour = 16'b00001_000001_00001; 
		1351: oled_colour = 16'b00001_000001_00001; 
		1352: oled_colour = 16'b00001_000001_00001; 
		1353: oled_colour = 16'b00001_000001_00001; 
		1354: oled_colour = 16'b00001_000001_00001; 
		1355: oled_colour = 16'b00001_000001_00001; 
		1356: oled_colour = 16'b00001_000001_00001; 
		1357: oled_colour = 16'b00001_000001_00001; 
		1358: oled_colour = 16'b00001_000001_00001; 
		1359: oled_colour = 16'b00001_000001_00001; 
		1360: oled_colour = 16'b00001_000001_00001; 
		1361: oled_colour = 16'b00001_000001_00001; 
		1362: oled_colour = 16'b00001_000001_00001; 
		1363: oled_colour = 16'b00001_000001_00001; 
		1364: oled_colour = 16'b00001_000001_00001; 
		1365: oled_colour = 16'b00001_000001_00001; 
		1366: oled_colour = 16'b00001_000001_00001; 
		1367: oled_colour = 16'b00001_000001_00001; 
		1368: oled_colour = 16'b00001_000001_00001; 
		1369: oled_colour = 16'b00001_000001_00001; 
		1370: oled_colour = 16'b00001_000001_00001; 
		1371: oled_colour = 16'b00001_000001_00001; 
		1372: oled_colour = 16'b00001_000001_00001; 
		1373: oled_colour = 16'b00001_000001_00001; 
		1374: oled_colour = 16'b00001_000001_00001; 
		1375: oled_colour = 16'b00001_000001_00001; 
		1376: oled_colour = 16'b00001_000001_00001; 
		1377: oled_colour = 16'b00001_000001_00001; 
		1378: oled_colour = 16'b00001_000001_00001; 
		1379: oled_colour = 16'b00001_000001_00001; 
		1380: oled_colour = 16'b00001_000001_00001; 
		1381: oled_colour = 16'b00001_000001_00001; 
		1382: oled_colour = 16'b00001_000001_00001; 
		1383: oled_colour = 16'b00001_000001_00001; 
		1384: oled_colour = 16'b00001_000001_00001; 
		1385: oled_colour = 16'b00001_000001_00001; 
		1386: oled_colour = 16'b00001_000001_00001; 
		1387: oled_colour = 16'b00001_000001_00001; 
		1388: oled_colour = 16'b00001_000001_00001; 
		1389: oled_colour = 16'b00001_000001_00001; 
		1390: oled_colour = 16'b00001_000001_00001; 
		1391: oled_colour = 16'b00001_000001_00001; 
		1392: oled_colour = 16'b00001_000001_00001; 
		1393: oled_colour = 16'b00001_000001_00001; 
		1394: oled_colour = 16'b00001_000001_00001; 
		1395: oled_colour = 16'b00001_000001_00001; 
		1396: oled_colour = 16'b00001_000001_00001; 
		1397: oled_colour = 16'b00001_000001_00001; 
		1398: oled_colour = 16'b00001_000001_00001; 
		1399: oled_colour = 16'b00001_000001_00001; 
		1400: oled_colour = 16'b00001_000001_00001; 
		1401: oled_colour = 16'b00001_000001_00001; 
		1402: oled_colour = 16'b00001_000001_00001; 
		1403: oled_colour = 16'b00001_000001_00001; 
		1404: oled_colour = 16'b00001_000001_00001; 
		1405: oled_colour = 16'b00001_000001_00001; 
		1406: oled_colour = 16'b00001_000001_00001; 
		1407: oled_colour = 16'b00001_000001_00001; 
		1408: oled_colour = 16'b00001_000001_00001; 
		1409: oled_colour = 16'b00001_000001_00001; 
		1410: oled_colour = 16'b00001_000001_00001; 
		1411: oled_colour = 16'b00001_000001_00001; 
		1412: oled_colour = 16'b00001_000001_00001; 
		1413: oled_colour = 16'b00001_000001_00001; 
		1414: oled_colour = 16'b00001_000001_00001; 
		1415: oled_colour = 16'b00001_000001_00001; 
		1416: oled_colour = 16'b00001_000001_00001; 
		1417: oled_colour = 16'b00001_000001_00001; 
		1418: oled_colour = 16'b00001_000001_00001; 
		1419: oled_colour = 16'b00001_000001_00001; 
		1420: oled_colour = 16'b00001_000001_00001; 
		1421: oled_colour = 16'b00001_000001_00001; 
		1422: oled_colour = 16'b00001_000001_00001; 
		1423: oled_colour = 16'b00001_000001_00001; 
		1424: oled_colour = 16'b00001_000001_00001; 
		1425: oled_colour = 16'b00001_000001_00001; 
		1426: oled_colour = 16'b00001_000001_00001; 
		1427: oled_colour = 16'b00001_000001_00001; 
		1428: oled_colour = 16'b00001_000001_00001; 
		1429: oled_colour = 16'b00001_000001_00001; 
		1430: oled_colour = 16'b00001_000001_00001; 
		1431: oled_colour = 16'b00001_000001_00001; 
		1432: oled_colour = 16'b00001_000001_00001; 
		1433: oled_colour = 16'b00001_000001_00001; 
		1434: oled_colour = 16'b00001_000001_00001; 
		1435: oled_colour = 16'b00001_000001_00001; 
		1436: oled_colour = 16'b00001_000001_00001; 
		1437: oled_colour = 16'b00001_000001_00001; 
		1438: oled_colour = 16'b00001_000001_00001; 
		1439: oled_colour = 16'b00001_000001_00001; 
		1440: oled_colour = 16'b00001_000001_00001; 
		1441: oled_colour = 16'b00001_000001_00001; 
		1442: oled_colour = 16'b00001_000001_00001; 
		1443: oled_colour = 16'b00001_000001_00001; 
		1444: oled_colour = 16'b00001_000001_00001; 
		1445: oled_colour = 16'b00001_000001_00001; 
		1446: oled_colour = 16'b00001_000001_00001; 
		1447: oled_colour = 16'b00001_000001_00001; 
		1448: oled_colour = 16'b00001_000001_00001; 
		1449: oled_colour = 16'b00001_000001_00001; 
		1450: oled_colour = 16'b00001_000001_00001; 
		1451: oled_colour = 16'b00001_000001_00001; 
		1452: oled_colour = 16'b00001_000001_00001; 
		1453: oled_colour = 16'b00001_000001_00001; 
		1454: oled_colour = 16'b00001_000001_00001; 
		1455: oled_colour = 16'b00001_000001_00001; 
		1456: oled_colour = 16'b00001_000001_00001; 
		1457: oled_colour = 16'b00001_000001_00001; 
		1458: oled_colour = 16'b00001_000001_00001; 
		1459: oled_colour = 16'b00001_000001_00001; 
		1460: oled_colour = 16'b00001_000001_00001; 
		1461: oled_colour = 16'b00001_000001_00001; 
		1462: oled_colour = 16'b00001_000001_00001; 
		1463: oled_colour = 16'b00001_000001_00001; 
		1464: oled_colour = 16'b00001_000001_00001; 
		1465: oled_colour = 16'b00001_000001_00001; 
		1466: oled_colour = 16'b00001_000001_00001; 
		1467: oled_colour = 16'b00001_000001_00001; 
		1468: oled_colour = 16'b00001_000001_00001; 
		1469: oled_colour = 16'b00001_000001_00001; 
		1470: oled_colour = 16'b00001_000001_00001; 
		1471: oled_colour = 16'b00001_000001_00001; 
		1472: oled_colour = 16'b00001_000001_00001; 
		1473: oled_colour = 16'b00001_000001_00001; 
		1474: oled_colour = 16'b11111_000001_00001; 
		1475: oled_colour = 16'b11111_111111_00001; 
		1476: oled_colour = 16'b11111_100000_10000; 
		1477: oled_colour = 16'b11000_100000_01000; 
		1478: oled_colour = 16'b11111_111111_01011; 
		1479: oled_colour = 16'b11000_110000_10000; 
		1480: oled_colour = 16'b11111_111111_11111; 
		1481: oled_colour = 16'b10110_111111_11111; 
		1482: oled_colour = 16'b11111_111111_11111; 
		1483: oled_colour = 16'b11111_111111_11111; 
		1484: oled_colour = 16'b11111_111111_11111; 
		1485: oled_colour = 16'b10110_111111_11111; 
		1486: oled_colour = 16'b10110_111111_11111; 
		1487: oled_colour = 16'b01011_101011_11111; 
		1488: oled_colour = 16'b10000_100000_11111; 
		1489: oled_colour = 16'b00001_111111_11111; 
		1490: oled_colour = 16'b00001_000001_11111; 
		1491: oled_colour = 16'b00001_000001_00001; 
		1492: oled_colour = 16'b00001_000001_00001; 
		1493: oled_colour = 16'b00001_000001_00001; 
		1494: oled_colour = 16'b00001_000001_00001; 
		1495: oled_colour = 16'b00001_000001_00001; 
		1496: oled_colour = 16'b00001_000001_00001; 
		1497: oled_colour = 16'b00001_000001_00001; 
		1498: oled_colour = 16'b00001_000001_00001; 
		1499: oled_colour = 16'b00001_000001_00001; 
		1500: oled_colour = 16'b00001_000001_00001; 
		1501: oled_colour = 16'b00001_000001_00001; 
		1502: oled_colour = 16'b00001_000001_00001; 
		1503: oled_colour = 16'b00001_000001_00001; 
		1504: oled_colour = 16'b00001_000001_00001; 
		1505: oled_colour = 16'b00001_000001_00001; 
		1506: oled_colour = 16'b00001_000001_00001; 
		1507: oled_colour = 16'b00001_000001_00001; 
		1508: oled_colour = 16'b00001_000001_00001; 
		1509: oled_colour = 16'b00001_000001_00001; 
		1510: oled_colour = 16'b00001_000001_00001; 
		1511: oled_colour = 16'b00001_000001_00001; 
		1512: oled_colour = 16'b00001_000001_00001; 
		1513: oled_colour = 16'b00001_000001_00001; 
		1514: oled_colour = 16'b00001_000001_00001; 
		1515: oled_colour = 16'b00001_000001_00001; 
		1516: oled_colour = 16'b00001_000001_00001; 
		1517: oled_colour = 16'b00001_000001_00001; 
		1518: oled_colour = 16'b00001_000001_00001; 
		1519: oled_colour = 16'b00001_000001_00001; 
		1520: oled_colour = 16'b00001_000001_00001; 
		1521: oled_colour = 16'b00001_000001_00001; 
		1522: oled_colour = 16'b00001_000001_00001; 
		1523: oled_colour = 16'b00001_000001_00001; 
		1524: oled_colour = 16'b00001_000001_00001; 
		1525: oled_colour = 16'b00001_000001_00001; 
		1526: oled_colour = 16'b00001_000001_00001; 
		1527: oled_colour = 16'b00001_000001_00001; 
		1528: oled_colour = 16'b00001_000001_00001; 
		1529: oled_colour = 16'b00001_000001_00001; 
		1530: oled_colour = 16'b00001_000001_00001; 
		1531: oled_colour = 16'b00001_000001_00001; 
		1532: oled_colour = 16'b00001_000001_00001; 
		1533: oled_colour = 16'b00001_000001_00001; 
		1534: oled_colour = 16'b00001_000001_00001; 
		1535: oled_colour = 16'b00001_000001_00001; 
		1536: oled_colour = 16'b00001_000001_00001; 
		1537: oled_colour = 16'b00001_000001_00001; 
		1538: oled_colour = 16'b00001_000001_00001; 
		1539: oled_colour = 16'b00001_000001_00001; 
		1540: oled_colour = 16'b00001_000001_00001; 
		1541: oled_colour = 16'b00001_000001_00001; 
		1542: oled_colour = 16'b00001_000001_00001; 
		1543: oled_colour = 16'b00001_000001_00001; 
		1544: oled_colour = 16'b00001_000001_00001; 
		1545: oled_colour = 16'b00001_000001_00001; 
		1546: oled_colour = 16'b00001_000001_00001; 
		1547: oled_colour = 16'b00001_000001_00001; 
		1548: oled_colour = 16'b00001_000001_00001; 
		1549: oled_colour = 16'b00001_000001_00001; 
		1550: oled_colour = 16'b00001_000001_00001; 
		1551: oled_colour = 16'b00001_000001_00001; 
		1552: oled_colour = 16'b00001_000001_00001; 
		1553: oled_colour = 16'b00001_000001_00001; 
		1554: oled_colour = 16'b00001_000001_00001; 
		1555: oled_colour = 16'b00001_000001_00001; 
		1556: oled_colour = 16'b00001_000001_00001; 
		1557: oled_colour = 16'b00001_000001_00001; 
		1558: oled_colour = 16'b00001_000001_00001; 
		1559: oled_colour = 16'b00001_000001_00001; 
		1560: oled_colour = 16'b00001_000001_00001; 
		1561: oled_colour = 16'b00001_000001_00001; 
		1562: oled_colour = 16'b00001_000001_00001; 
		1563: oled_colour = 16'b00001_000001_00001; 
		1564: oled_colour = 16'b00001_000001_00001; 
		1565: oled_colour = 16'b00001_000001_00001; 
		1566: oled_colour = 16'b00001_000001_00001; 
		1567: oled_colour = 16'b00001_000001_00001; 
		1568: oled_colour = 16'b00001_000001_00001; 
		1569: oled_colour = 16'b00001_000001_00001; 
		1570: oled_colour = 16'b00001_000001_00001; 
		1571: oled_colour = 16'b00001_000001_00001; 
		1572: oled_colour = 16'b00001_000001_00001; 
		1573: oled_colour = 16'b00001_000001_00001; 
		1574: oled_colour = 16'b00001_000001_00001; 
		1575: oled_colour = 16'b00001_000001_00001; 
		1576: oled_colour = 16'b00001_000001_00001; 
		1577: oled_colour = 16'b00001_000001_00001; 
		1578: oled_colour = 16'b00001_000001_00001; 
		1579: oled_colour = 16'b00001_000001_00001; 
		1580: oled_colour = 16'b00001_000001_00001; 
		1581: oled_colour = 16'b00001_000001_00001; 
		1582: oled_colour = 16'b00001_000001_00001; 
		1583: oled_colour = 16'b00001_000001_00001; 
		1584: oled_colour = 16'b00001_000001_00001; 
		1585: oled_colour = 16'b00001_000001_00001; 
		1586: oled_colour = 16'b00001_000001_00001; 
		1587: oled_colour = 16'b11111_111111_11111; 
		1588: oled_colour = 16'b01000_100000_11000; 
		1589: oled_colour = 16'b01011_101011_11111; 
		1590: oled_colour = 16'b00001_100000_10000; 
		1591: oled_colour = 16'b00001_000001_00001; 
		1592: oled_colour = 16'b00001_000001_00001; 
		1593: oled_colour = 16'b00001_000001_00001; 
		1594: oled_colour = 16'b00001_000001_00001; 
		1595: oled_colour = 16'b00001_000001_00001; 
		1596: oled_colour = 16'b00001_000001_00001; 
		1597: oled_colour = 16'b00001_000001_00001; 
		1598: oled_colour = 16'b00001_000001_00001; 
		1599: oled_colour = 16'b00001_000001_00001; 
		1600: oled_colour = 16'b00001_000001_00001; 
		1601: oled_colour = 16'b00001_000001_00001; 
		1602: oled_colour = 16'b00001_000001_00001; 
		1603: oled_colour = 16'b00001_000001_00001; 
		1604: oled_colour = 16'b00001_000001_00001; 
		1605: oled_colour = 16'b00001_000001_00001; 
		1606: oled_colour = 16'b00001_000001_00001; 
		1607: oled_colour = 16'b00001_000001_00001; 
		1608: oled_colour = 16'b00001_000001_00001; 
		1609: oled_colour = 16'b00001_000001_00001; 
		1610: oled_colour = 16'b00001_000001_00001; 
		1611: oled_colour = 16'b00001_000001_00001; 
		1612: oled_colour = 16'b00001_000001_00001; 
		1613: oled_colour = 16'b00001_000001_00001; 
		1614: oled_colour = 16'b00001_000001_00001; 
		1615: oled_colour = 16'b00001_000001_00001; 
		1616: oled_colour = 16'b00001_000001_00001; 
		1617: oled_colour = 16'b00001_000001_00001; 
		1618: oled_colour = 16'b00001_000001_00001; 
		1619: oled_colour = 16'b00001_000001_00001; 
		1620: oled_colour = 16'b00001_000001_00001; 
		1621: oled_colour = 16'b00001_000001_00001; 
		1622: oled_colour = 16'b00001_000001_00001; 
		1623: oled_colour = 16'b00001_000001_00001; 
		1624: oled_colour = 16'b00001_000001_00001; 
		1625: oled_colour = 16'b00001_000001_00001; 
		1626: oled_colour = 16'b00001_000001_00001; 
		1627: oled_colour = 16'b00001_000001_00001; 
		1628: oled_colour = 16'b00001_000001_00001; 
		1629: oled_colour = 16'b00001_000001_00001; 
		1630: oled_colour = 16'b00001_000001_00001; 
		1631: oled_colour = 16'b00001_000001_00001; 
		1632: oled_colour = 16'b00001_000001_00001; 
		1633: oled_colour = 16'b00001_000001_00001; 
		1634: oled_colour = 16'b00001_000001_00001; 
		1635: oled_colour = 16'b00001_000001_00001; 
		1636: oled_colour = 16'b00001_000001_00001; 
		1637: oled_colour = 16'b00001_000001_00001; 
		1638: oled_colour = 16'b00001_000001_00001; 
		1639: oled_colour = 16'b00001_000001_00001; 
		1640: oled_colour = 16'b00001_000001_00001; 
		1641: oled_colour = 16'b00001_000001_00001; 
		1642: oled_colour = 16'b00001_000001_00001; 
		1643: oled_colour = 16'b00001_000001_00001; 
		1644: oled_colour = 16'b00001_000001_00001; 
		1645: oled_colour = 16'b00001_000001_00001; 
		1646: oled_colour = 16'b00001_000001_00001; 
		1647: oled_colour = 16'b00001_000001_00001; 
		1648: oled_colour = 16'b00001_000001_00001; 
		1649: oled_colour = 16'b00001_000001_00001; 
		1650: oled_colour = 16'b00001_000001_00001; 
		1651: oled_colour = 16'b00001_000001_00001; 
		1652: oled_colour = 16'b00001_000001_00001; 
		1653: oled_colour = 16'b00001_000001_00001; 
		1654: oled_colour = 16'b00001_000001_00001; 
		1655: oled_colour = 16'b00001_000001_00001; 
		1656: oled_colour = 16'b00001_000001_00001; 
		1657: oled_colour = 16'b00001_000001_00001; 
		1658: oled_colour = 16'b00001_000001_00001; 
		1659: oled_colour = 16'b00001_000001_00001; 
		1660: oled_colour = 16'b00001_000001_00001; 
		1661: oled_colour = 16'b00001_000001_00001; 
		1662: oled_colour = 16'b00001_000001_00001; 
		1663: oled_colour = 16'b00001_000001_00001; 
		1664: oled_colour = 16'b00001_000001_00001; 
		1665: oled_colour = 16'b10110_010110_01011; 
		1666: oled_colour = 16'b11000_011101_01010; 
		1667: oled_colour = 16'b10111_101001_01101; 
		1668: oled_colour = 16'b11001_100010_01100; 
		1669: oled_colour = 16'b11011_100101_01100; 
		1670: oled_colour = 16'b11010_101111_01111; 
		1671: oled_colour = 16'b11011_110110_10101; 
		1672: oled_colour = 16'b11010_110101_11011; 
		1673: oled_colour = 16'b11000_110110_11111; 
		1674: oled_colour = 16'b10111_111000_11111; 
		1675: oled_colour = 16'b10111_110111_11111; 
		1676: oled_colour = 16'b10111_110110_11111; 
		1677: oled_colour = 16'b10100_110010_11111; 
		1678: oled_colour = 16'b10000_101100_11110; 
		1679: oled_colour = 16'b01100_100110_11011; 
		1680: oled_colour = 16'b00101_011110_11001; 
		1681: oled_colour = 16'b00001_000101_10101; 
		1682: oled_colour = 16'b00001_000001_00001; 
		1683: oled_colour = 16'b00001_000001_00001; 
		1684: oled_colour = 16'b00001_000001_00001; 
		1685: oled_colour = 16'b00001_000001_00001; 
		1686: oled_colour = 16'b00001_000001_00001; 
		1687: oled_colour = 16'b00001_100000_11111; 
		1688: oled_colour = 16'b00001_010110_10110; 
		1689: oled_colour = 16'b00001_000001_00001; 
		1690: oled_colour = 16'b00001_000001_00001; 
		1691: oled_colour = 16'b00001_000001_00001; 
		1692: oled_colour = 16'b00001_000001_00001; 
		1693: oled_colour = 16'b00001_000001_00001; 
		1694: oled_colour = 16'b00001_000001_00001; 
		1695: oled_colour = 16'b00001_000001_00001; 
		1696: oled_colour = 16'b00001_000001_00001; 
		1697: oled_colour = 16'b00001_000001_00001; 
		1698: oled_colour = 16'b00001_000001_00001; 
		1699: oled_colour = 16'b00001_000001_00001; 
		1700: oled_colour = 16'b00001_000001_00001; 
		1701: oled_colour = 16'b00001_000001_00001; 
		1702: oled_colour = 16'b00001_000001_00001; 
		1703: oled_colour = 16'b00001_000001_00001; 
		1704: oled_colour = 16'b00001_000001_00001; 
		1705: oled_colour = 16'b00001_000001_00001; 
		1706: oled_colour = 16'b00001_000001_00001; 
		1707: oled_colour = 16'b00001_000001_00001; 
		1708: oled_colour = 16'b00001_000001_00001; 
		1709: oled_colour = 16'b00001_000001_00001; 
		1710: oled_colour = 16'b00001_000001_00001; 
		1711: oled_colour = 16'b00001_000001_00001; 
		1712: oled_colour = 16'b00001_000001_00001; 
		1713: oled_colour = 16'b00001_000001_00001; 
		1714: oled_colour = 16'b00001_000001_00001; 
		1715: oled_colour = 16'b00001_000001_00001; 
		1716: oled_colour = 16'b00001_000001_00001; 
		1717: oled_colour = 16'b00001_000001_00001; 
		1718: oled_colour = 16'b00001_000001_00001; 
		1719: oled_colour = 16'b00001_000001_00001; 
		1720: oled_colour = 16'b00001_000001_00001; 
		1721: oled_colour = 16'b00001_000001_00001; 
		1722: oled_colour = 16'b00001_000001_00001; 
		1723: oled_colour = 16'b00001_000001_00001; 
		1724: oled_colour = 16'b00001_000001_00001; 
		1725: oled_colour = 16'b00001_000001_00001; 
		1726: oled_colour = 16'b00001_000001_00001; 
		1727: oled_colour = 16'b00001_000001_00001; 
		1728: oled_colour = 16'b00001_000001_00001; 
		1729: oled_colour = 16'b00001_000001_00001; 
		1730: oled_colour = 16'b00001_000001_00001; 
		1731: oled_colour = 16'b00001_000001_00001; 
		1732: oled_colour = 16'b00001_000001_00001; 
		1733: oled_colour = 16'b00001_000001_00001; 
		1734: oled_colour = 16'b00001_000001_00001; 
		1735: oled_colour = 16'b00001_000001_00001; 
		1736: oled_colour = 16'b00001_000001_00001; 
		1737: oled_colour = 16'b00001_000001_00001; 
		1738: oled_colour = 16'b00001_000001_00001; 
		1739: oled_colour = 16'b00001_000001_00001; 
		1740: oled_colour = 16'b00001_000001_00001; 
		1741: oled_colour = 16'b00001_000001_00001; 
		1742: oled_colour = 16'b00001_000001_00001; 
		1743: oled_colour = 16'b00001_000001_00001; 
		1744: oled_colour = 16'b00001_000001_00001; 
		1745: oled_colour = 16'b00001_000001_00001; 
		1746: oled_colour = 16'b00001_000001_00001; 
		1747: oled_colour = 16'b00001_000001_00001; 
		1748: oled_colour = 16'b00001_000001_00001; 
		1749: oled_colour = 16'b00001_000001_00001; 
		1750: oled_colour = 16'b00001_000001_00001; 
		1751: oled_colour = 16'b00001_000001_00001; 
		1752: oled_colour = 16'b00001_000001_00001; 
		1753: oled_colour = 16'b00001_000001_00001; 
		1754: oled_colour = 16'b00001_000001_00001; 
		1755: oled_colour = 16'b00001_000001_00001; 
		1756: oled_colour = 16'b00001_000001_00001; 
		1757: oled_colour = 16'b00001_000001_00001; 
		1758: oled_colour = 16'b00001_000001_00001; 
		1759: oled_colour = 16'b00001_000001_00001; 
		1760: oled_colour = 16'b00001_000001_11111; 
		1761: oled_colour = 16'b10110_010100_01010; 
		1762: oled_colour = 16'b11000_011110_01000; 
		1763: oled_colour = 16'b11000_101011_01100; 
		1764: oled_colour = 16'b11010_100111_01100; 
		1765: oled_colour = 16'b11101_101010_01101; 
		1766: oled_colour = 16'b11101_110010_10000; 
		1767: oled_colour = 16'b11101_111000_10100; 
		1768: oled_colour = 16'b11100_111001_10110; 
		1769: oled_colour = 16'b11100_111001_11001; 
		1770: oled_colour = 16'b11101_111000_11000; 
		1771: oled_colour = 16'b11111_111100_11010; 
		1772: oled_colour = 16'b11111_111111_11011; 
		1773: oled_colour = 16'b11111_111111_11110; 
		1774: oled_colour = 16'b11110_111111_11111; 
		1775: oled_colour = 16'b11010_111100_11111; 
		1776: oled_colour = 16'b10111_110110_11111; 
		1777: oled_colour = 16'b10101_110100_11110; 
		1778: oled_colour = 16'b10000_101111_11101; 
		1779: oled_colour = 16'b01100_101001_11100; 
		1780: oled_colour = 16'b01001_100010_11011; 
		1781: oled_colour = 16'b00110_011011_11001; 
		1782: oled_colour = 16'b00100_010010_10110; 
		1783: oled_colour = 16'b00001_000001_00001; 
		1784: oled_colour = 16'b00001_000001_00001; 
		1785: oled_colour = 16'b00001_100000_10000; 
		1786: oled_colour = 16'b00001_000001_00001; 
		1787: oled_colour = 16'b00001_000001_00001; 
		1788: oled_colour = 16'b00001_000001_00001; 
		1789: oled_colour = 16'b00001_000001_00001; 
		1790: oled_colour = 16'b00001_000001_00001; 
		1791: oled_colour = 16'b00001_000001_00001; 
		1792: oled_colour = 16'b00001_000001_00001; 
		1793: oled_colour = 16'b00001_000001_00001; 
		1794: oled_colour = 16'b00001_000001_00001; 
		1795: oled_colour = 16'b00001_000001_00001; 
		1796: oled_colour = 16'b00001_000001_00001; 
		1797: oled_colour = 16'b00001_000001_00001; 
		1798: oled_colour = 16'b00001_000001_00001; 
		1799: oled_colour = 16'b00001_000001_00001; 
		1800: oled_colour = 16'b00001_000001_00001; 
		1801: oled_colour = 16'b00001_000001_00001; 
		1802: oled_colour = 16'b00001_000001_00001; 
		1803: oled_colour = 16'b00001_000001_00001; 
		1804: oled_colour = 16'b00001_000001_00001; 
		1805: oled_colour = 16'b00001_000001_00001; 
		1806: oled_colour = 16'b00001_000001_00001; 
		1807: oled_colour = 16'b00001_000001_00001; 
		1808: oled_colour = 16'b00001_000001_00001; 
		1809: oled_colour = 16'b00001_000001_00001; 
		1810: oled_colour = 16'b00001_000001_00001; 
		1811: oled_colour = 16'b00001_000001_00001; 
		1812: oled_colour = 16'b00001_000001_00001; 
		1813: oled_colour = 16'b00001_000001_00001; 
		1814: oled_colour = 16'b00001_000001_00001; 
		1815: oled_colour = 16'b00001_000001_00001; 
		1816: oled_colour = 16'b00001_000001_00001; 
		1817: oled_colour = 16'b00001_000001_00001; 
		1818: oled_colour = 16'b00001_000001_00001; 
		1819: oled_colour = 16'b00001_000001_00001; 
		1820: oled_colour = 16'b00001_000001_00001; 
		1821: oled_colour = 16'b00001_000001_00001; 
		1822: oled_colour = 16'b00001_000001_00001; 
		1823: oled_colour = 16'b00001_000001_00001; 
		1824: oled_colour = 16'b00001_000001_00001; 
		1825: oled_colour = 16'b00001_000001_00001; 
		1826: oled_colour = 16'b00001_000001_00001; 
		1827: oled_colour = 16'b00001_000001_00001; 
		1828: oled_colour = 16'b00001_000001_00001; 
		1829: oled_colour = 16'b00001_000001_00001; 
		1830: oled_colour = 16'b00001_000001_00001; 
		1831: oled_colour = 16'b00001_000001_00001; 
		1832: oled_colour = 16'b00001_000001_00001; 
		1833: oled_colour = 16'b00001_000001_00001; 
		1834: oled_colour = 16'b00001_000001_00001; 
		1835: oled_colour = 16'b00001_000001_00001; 
		1836: oled_colour = 16'b00001_000001_00001; 
		1837: oled_colour = 16'b00001_000001_00001; 
		1838: oled_colour = 16'b00001_000001_00001; 
		1839: oled_colour = 16'b00001_000001_00001; 
		1840: oled_colour = 16'b00001_000001_00001; 
		1841: oled_colour = 16'b00001_000001_00001; 
		1842: oled_colour = 16'b00001_000001_00001; 
		1843: oled_colour = 16'b00001_000001_00001; 
		1844: oled_colour = 16'b00001_000001_00001; 
		1845: oled_colour = 16'b00001_000001_00001; 
		1846: oled_colour = 16'b00001_000001_00001; 
		1847: oled_colour = 16'b00001_000001_00001; 
		1848: oled_colour = 16'b00001_000001_00001; 
		1849: oled_colour = 16'b00001_000001_00001; 
		1850: oled_colour = 16'b00001_000001_00001; 
		1851: oled_colour = 16'b00001_000001_00001; 
		1852: oled_colour = 16'b00001_000001_00001; 
		1853: oled_colour = 16'b00001_000001_00001; 
		1854: oled_colour = 16'b00001_000001_00001; 
		1855: oled_colour = 16'b00001_000001_00001; 
		1856: oled_colour = 16'b00001_000001_00001; 
		1857: oled_colour = 16'b00001_000001_00001; 
		1858: oled_colour = 16'b00001_000001_00001; 
		1859: oled_colour = 16'b00001_000001_00001; 
		1860: oled_colour = 16'b00001_000001_00001; 
		1861: oled_colour = 16'b00001_000001_00001; 
		1862: oled_colour = 16'b00001_000001_00001; 
		1863: oled_colour = 16'b00001_000001_00001; 
		1864: oled_colour = 16'b01010_001010_00001; 
		1865: oled_colour = 16'b01000_000001_00001; 
		1866: oled_colour = 16'b10111_010101_00110; 
		1867: oled_colour = 16'b11010_011111_00110; 
		1868: oled_colour = 16'b11010_100111_01001; 
		1869: oled_colour = 16'b11100_101001_01011; 
		1870: oled_colour = 16'b11101_101100_01100; 
		1871: oled_colour = 16'b11111_110110_01111; 
		1872: oled_colour = 16'b11111_111110_10100; 
		1873: oled_colour = 16'b11111_111111_11100; 
		1874: oled_colour = 16'b11110_111111_11111; 
		1875: oled_colour = 16'b11010_111101_11111; 
		1876: oled_colour = 16'b10100_111000_11111; 
		1877: oled_colour = 16'b01110_101110_11110; 
		1878: oled_colour = 16'b01001_100010_11011; 
		1879: oled_colour = 16'b00110_011011_11001; 
		1880: oled_colour = 16'b00100_010010_10110; 
		1881: oled_colour = 16'b00001_000001_00001; 
		1882: oled_colour = 16'b00001_000001_00001; 
		1883: oled_colour = 16'b00001_000001_00001; 
		1884: oled_colour = 16'b00001_000001_00001; 
		1885: oled_colour = 16'b00001_000001_00001; 
		1886: oled_colour = 16'b00001_000001_00001; 
		1887: oled_colour = 16'b00001_000001_00001; 
		1888: oled_colour = 16'b00001_000001_00001; 
		1889: oled_colour = 16'b00001_000001_00001; 
		1890: oled_colour = 16'b00001_000001_00001; 
		1891: oled_colour = 16'b00001_000001_00001; 
		1892: oled_colour = 16'b00001_000001_00001; 
		1893: oled_colour = 16'b00001_000001_00001; 
		1894: oled_colour = 16'b00001_000001_00001; 
		1895: oled_colour = 16'b00001_000001_00001; 
		1896: oled_colour = 16'b00001_000001_00001; 
		1897: oled_colour = 16'b00001_000001_00001; 
		1898: oled_colour = 16'b00001_000001_00001; 
		1899: oled_colour = 16'b00001_000001_00001; 
		1900: oled_colour = 16'b00001_000001_00001; 
		1901: oled_colour = 16'b00001_000001_00001; 
		1902: oled_colour = 16'b00001_000001_00001; 
		1903: oled_colour = 16'b00001_000001_00001; 
		1904: oled_colour = 16'b00001_000001_00001; 
		1905: oled_colour = 16'b00001_000001_00001; 
		1906: oled_colour = 16'b00001_000001_00001; 
		1907: oled_colour = 16'b00001_000001_00001; 
		1908: oled_colour = 16'b00001_000001_00001; 
		1909: oled_colour = 16'b00001_000001_00001; 
		1910: oled_colour = 16'b00001_000001_00001; 
		1911: oled_colour = 16'b00001_000001_00001; 
		1912: oled_colour = 16'b00001_000001_00001; 
		1913: oled_colour = 16'b00001_000001_00001; 
		1914: oled_colour = 16'b00001_000001_00001; 
		1915: oled_colour = 16'b00001_000001_00001; 
		1916: oled_colour = 16'b00001_000001_00001; 
		1917: oled_colour = 16'b00001_000001_00001; 
		1918: oled_colour = 16'b00001_000001_00001; 
		1919: oled_colour = 16'b00001_000001_00001; 
		1920: oled_colour = 16'b00001_000001_00001; 
		1921: oled_colour = 16'b00001_000001_00001; 
		1922: oled_colour = 16'b00001_000001_00001; 
		1923: oled_colour = 16'b00001_000001_00001; 
		1924: oled_colour = 16'b00001_000001_00001; 
		1925: oled_colour = 16'b00001_000001_00001; 
		1926: oled_colour = 16'b00001_000001_00001; 
		1927: oled_colour = 16'b00001_000001_00001; 
		1928: oled_colour = 16'b00001_000001_00001; 
		1929: oled_colour = 16'b00001_000001_00001; 
		1930: oled_colour = 16'b00001_000001_00001; 
		1931: oled_colour = 16'b00001_000001_00001; 
		1932: oled_colour = 16'b00001_000001_00001; 
		1933: oled_colour = 16'b00001_000001_00001; 
		1934: oled_colour = 16'b00001_000001_00001; 
		1935: oled_colour = 16'b00001_000001_00001; 
		1936: oled_colour = 16'b00001_000001_00001; 
		1937: oled_colour = 16'b00001_000001_00001; 
		1938: oled_colour = 16'b00001_000001_00001; 
		1939: oled_colour = 16'b00001_000001_00001; 
		1940: oled_colour = 16'b00001_000001_00001; 
		1941: oled_colour = 16'b00001_000001_00001; 
		1942: oled_colour = 16'b00001_000001_00001; 
		1943: oled_colour = 16'b00001_000001_00001; 
		1944: oled_colour = 16'b00001_000001_00001; 
		1945: oled_colour = 16'b00001_000001_00001; 
		1946: oled_colour = 16'b00001_000001_00001; 
		1947: oled_colour = 16'b00001_000001_00001; 
		1948: oled_colour = 16'b00001_000001_00001; 
		1949: oled_colour = 16'b00001_000001_00001; 
		1950: oled_colour = 16'b00001_000001_00001; 
		1951: oled_colour = 16'b00001_000001_00001; 
		1952: oled_colour = 16'b00001_000001_00001; 
		1953: oled_colour = 16'b10000_100000_00001; 
		1954: oled_colour = 16'b11111_100000_00001; 
		1955: oled_colour = 16'b11111_100000_10000; 
		1956: oled_colour = 16'b00001_000001_00001; 
		1957: oled_colour = 16'b00001_000001_00001; 
		1958: oled_colour = 16'b00001_000001_00001; 
		1959: oled_colour = 16'b00001_000001_00001; 
		1960: oled_colour = 16'b00001_000001_00001; 
		1961: oled_colour = 16'b00001_000001_00001; 
		1962: oled_colour = 16'b00001_000001_00001; 
		1963: oled_colour = 16'b00001_000001_00001; 
		1964: oled_colour = 16'b00001_000001_00001; 
		1965: oled_colour = 16'b00001_000001_00001; 
		1966: oled_colour = 16'b01111_000001_00001; 
		1967: oled_colour = 16'b11010_011010_00011; 
		1968: oled_colour = 16'b11101_101010_00101; 
		1969: oled_colour = 16'b11111_111011_01110; 
		1970: oled_colour = 16'b11111_111101_11001; 
		1971: oled_colour = 16'b11111_111101_11110; 
		1972: oled_colour = 16'b11110_111110_11111; 
		1973: oled_colour = 16'b11010_111100_11111; 
		1974: oled_colour = 16'b10100_110111_11111; 
		1975: oled_colour = 16'b01111_101111_11111; 
		1976: oled_colour = 16'b01011_100110_11100; 
		1977: oled_colour = 16'b00111_011101_11001; 
		1978: oled_colour = 16'b00100_001101_10100; 
		1979: oled_colour = 16'b00001_000001_11111; 
		1980: oled_colour = 16'b00001_000001_00001; 
		1981: oled_colour = 16'b00001_000001_00001; 
		1982: oled_colour = 16'b00001_000001_00001; 
		1983: oled_colour = 16'b00001_000001_00001; 
		1984: oled_colour = 16'b00001_000001_00001; 
		1985: oled_colour = 16'b00001_000001_00001; 
		1986: oled_colour = 16'b00001_000001_00001; 
		1987: oled_colour = 16'b00001_000001_00001; 
		1988: oled_colour = 16'b00001_000001_00001; 
		1989: oled_colour = 16'b00001_000001_00001; 
		1990: oled_colour = 16'b00001_000001_00001; 
		1991: oled_colour = 16'b00001_000001_00001; 
		1992: oled_colour = 16'b00001_000001_00001; 
		1993: oled_colour = 16'b00001_000001_00001; 
		1994: oled_colour = 16'b00001_000001_00001; 
		1995: oled_colour = 16'b00001_000001_00001; 
		1996: oled_colour = 16'b00001_000001_00001; 
		1997: oled_colour = 16'b00001_000001_00001; 
		1998: oled_colour = 16'b00001_000001_00001; 
		1999: oled_colour = 16'b00001_000001_00001; 
		2000: oled_colour = 16'b00001_000001_00001; 
		2001: oled_colour = 16'b00001_000001_00001; 
		2002: oled_colour = 16'b00001_000001_00001; 
		2003: oled_colour = 16'b00001_000001_00001; 
		2004: oled_colour = 16'b00001_000001_00001; 
		2005: oled_colour = 16'b00001_000001_00001; 
		2006: oled_colour = 16'b00001_000001_00001; 
		2007: oled_colour = 16'b00001_000001_00001; 
		2008: oled_colour = 16'b00001_000001_00001; 
		2009: oled_colour = 16'b00001_000001_00001; 
		2010: oled_colour = 16'b00001_000001_00001; 
		2011: oled_colour = 16'b00001_000001_00001; 
		2012: oled_colour = 16'b00001_000001_00001; 
		2013: oled_colour = 16'b00001_000001_00001; 
		2014: oled_colour = 16'b00001_000001_00001; 
		2015: oled_colour = 16'b00001_000001_00001; 
		2016: oled_colour = 16'b00001_000001_00001; 
		2017: oled_colour = 16'b00001_000001_00001; 
		2018: oled_colour = 16'b00001_000001_00001; 
		2019: oled_colour = 16'b00001_000001_00001; 
		2020: oled_colour = 16'b00001_000001_00001; 
		2021: oled_colour = 16'b00001_000001_00001; 
		2022: oled_colour = 16'b00001_000001_00001; 
		2023: oled_colour = 16'b00001_000001_00001; 
		2024: oled_colour = 16'b00001_000001_00001; 
		2025: oled_colour = 16'b00001_000001_00001; 
		2026: oled_colour = 16'b00001_000001_00001; 
		2027: oled_colour = 16'b00001_000001_00001; 
		2028: oled_colour = 16'b00001_000001_00001; 
		2029: oled_colour = 16'b00001_000001_00001; 
		2030: oled_colour = 16'b00001_000001_00001; 
		2031: oled_colour = 16'b00001_000001_00001; 
		2032: oled_colour = 16'b00001_000001_00001; 
		2033: oled_colour = 16'b00001_000001_00001; 
		2034: oled_colour = 16'b00001_000001_00001; 
		2035: oled_colour = 16'b00001_000001_00001; 
		2036: oled_colour = 16'b00001_000001_00001; 
		2037: oled_colour = 16'b00001_000001_00001; 
		2038: oled_colour = 16'b00001_000001_00001; 
		2039: oled_colour = 16'b00001_000001_00001; 
		2040: oled_colour = 16'b00001_000001_00001; 
		2041: oled_colour = 16'b00001_000001_00001; 
		2042: oled_colour = 16'b00001_000001_00001; 
		2043: oled_colour = 16'b00001_000001_00001; 
		2044: oled_colour = 16'b00001_000001_00001; 
		2045: oled_colour = 16'b00001_000001_00001; 
		2046: oled_colour = 16'b00001_000001_00001; 
		2047: oled_colour = 16'b00001_000001_00001; 
		2048: oled_colour = 16'b00001_000001_00001; 
		2049: oled_colour = 16'b00001_000001_00001; 
		2050: oled_colour = 16'b00001_000001_00001; 
		2051: oled_colour = 16'b00001_000001_00001; 
		2052: oled_colour = 16'b00001_000001_00001; 
		2053: oled_colour = 16'b11111_000001_00001; 
		2054: oled_colour = 16'b11111_000001_00001; 
		2055: oled_colour = 16'b11111_111111_00001; 
		2056: oled_colour = 16'b11111_111111_00001; 
		2057: oled_colour = 16'b11111_111111_00001; 
		2058: oled_colour = 16'b11111_100000_10000; 
		2059: oled_colour = 16'b11111_101011_01011; 
		2060: oled_colour = 16'b11111_101011_01011; 
		2061: oled_colour = 16'b11111_111111_01011; 
		2062: oled_colour = 16'b00001_000001_00001; 
		2063: oled_colour = 16'b00001_000001_00001; 
		2064: oled_colour = 16'b11000_010100_00110; 
		2065: oled_colour = 16'b11111_110100_01001; 
		2066: oled_colour = 16'b11110_111110_10111; 
		2067: oled_colour = 16'b11110_111100_11110; 
		2068: oled_colour = 16'b11111_111101_11111; 
		2069: oled_colour = 16'b11111_111101_11110; 
		2070: oled_colour = 16'b11101_111101_11111; 
		2071: oled_colour = 16'b10111_111011_11111; 
		2072: oled_colour = 16'b10010_110101_11111; 
		2073: oled_colour = 16'b01010_100110_11101; 
		2074: oled_colour = 16'b00100_010100_10111; 
		2075: oled_colour = 16'b00001_000001_00001; 
		2076: oled_colour = 16'b00001_010110_10110; 
		2077: oled_colour = 16'b00001_000001_00001; 
		2078: oled_colour = 16'b00001_000001_00001; 
		2079: oled_colour = 16'b00001_000001_00001; 
		2080: oled_colour = 16'b00001_000001_00001; 
		2081: oled_colour = 16'b00001_000001_00001; 
		2082: oled_colour = 16'b00001_000001_00001; 
		2083: oled_colour = 16'b00001_000001_00001; 
		2084: oled_colour = 16'b00001_000001_00001; 
		2085: oled_colour = 16'b00001_000001_00001; 
		2086: oled_colour = 16'b00001_000001_00001; 
		2087: oled_colour = 16'b00001_000001_00001; 
		2088: oled_colour = 16'b00001_000001_00001; 
		2089: oled_colour = 16'b00001_000001_00001; 
		2090: oled_colour = 16'b00001_000001_00001; 
		2091: oled_colour = 16'b00001_000001_00001; 
		2092: oled_colour = 16'b00001_000001_00001; 
		2093: oled_colour = 16'b00001_000001_00001; 
		2094: oled_colour = 16'b00001_000001_00001; 
		2095: oled_colour = 16'b00001_000001_00001; 
		2096: oled_colour = 16'b00001_000001_00001; 
		2097: oled_colour = 16'b00001_000001_00001; 
		2098: oled_colour = 16'b00001_000001_00001; 
		2099: oled_colour = 16'b00001_000001_00001; 
		2100: oled_colour = 16'b00001_000001_00001; 
		2101: oled_colour = 16'b00001_000001_00001; 
		2102: oled_colour = 16'b00001_000001_00001; 
		2103: oled_colour = 16'b00001_000001_00001; 
		2104: oled_colour = 16'b00001_000001_00001; 
		2105: oled_colour = 16'b00001_000001_00001; 
		2106: oled_colour = 16'b00001_000001_00001; 
		2107: oled_colour = 16'b00001_000001_00001; 
		2108: oled_colour = 16'b00001_000001_00001; 
		2109: oled_colour = 16'b00001_000001_00001; 
		2110: oled_colour = 16'b00001_000001_00001; 
		2111: oled_colour = 16'b00001_000001_00001; 
		2112: oled_colour = 16'b00001_000001_00001; 
		2113: oled_colour = 16'b00001_000001_00001; 
		2114: oled_colour = 16'b00001_000001_00001; 
		2115: oled_colour = 16'b00001_000001_00001; 
		2116: oled_colour = 16'b00001_000001_00001; 
		2117: oled_colour = 16'b00001_000001_00001; 
		2118: oled_colour = 16'b00001_000001_00001; 
		2119: oled_colour = 16'b00001_000001_00001; 
		2120: oled_colour = 16'b00001_000001_00001; 
		2121: oled_colour = 16'b00001_000001_00001; 
		2122: oled_colour = 16'b00001_000001_00001; 
		2123: oled_colour = 16'b00001_000001_00001; 
		2124: oled_colour = 16'b00001_000001_00001; 
		2125: oled_colour = 16'b00001_000001_00001; 
		2126: oled_colour = 16'b00001_000001_00001; 
		2127: oled_colour = 16'b00001_000001_00001; 
		2128: oled_colour = 16'b00001_000001_00001; 
		2129: oled_colour = 16'b00001_000001_00001; 
		2130: oled_colour = 16'b00001_000001_00001; 
		2131: oled_colour = 16'b00001_000001_00001; 
		2132: oled_colour = 16'b00001_000001_00001; 
		2133: oled_colour = 16'b00001_000001_00001; 
		2134: oled_colour = 16'b00001_000001_00001; 
		2135: oled_colour = 16'b00001_000001_00001; 
		2136: oled_colour = 16'b00001_000001_00001; 
		2137: oled_colour = 16'b00001_000001_00001; 
		2138: oled_colour = 16'b00001_000001_00001; 
		2139: oled_colour = 16'b00001_000001_00001; 
		2140: oled_colour = 16'b00001_000001_00001; 
		2141: oled_colour = 16'b00001_000001_00001; 
		2142: oled_colour = 16'b00001_000001_00001; 
		2143: oled_colour = 16'b00001_000001_00001; 
		2144: oled_colour = 16'b00001_000001_00001; 
		2145: oled_colour = 16'b00001_000001_00001; 
		2146: oled_colour = 16'b00001_000001_00001; 
		2147: oled_colour = 16'b00001_000001_00001; 
		2148: oled_colour = 16'b00001_000001_00001; 
		2149: oled_colour = 16'b00001_000001_00001; 
		2150: oled_colour = 16'b00001_000001_00001; 
		2151: oled_colour = 16'b00001_000001_00001; 
		2152: oled_colour = 16'b00001_000001_00001; 
		2153: oled_colour = 16'b00001_000001_00001; 
		2154: oled_colour = 16'b00001_000001_00001; 
		2155: oled_colour = 16'b00001_000001_00001; 
		2156: oled_colour = 16'b00001_000001_00001; 
		2157: oled_colour = 16'b11111_100000_00001; 
		2158: oled_colour = 16'b10000_000001_11111; 
		2159: oled_colour = 16'b11001_011000_00111; 
		2160: oled_colour = 16'b11110_101010_00110; 
		2161: oled_colour = 16'b11111_111100_10000; 
		2162: oled_colour = 16'b11110_111100_11011; 
		2163: oled_colour = 16'b11110_111100_11111; 
		2164: oled_colour = 16'b11111_111100_11110; 
		2165: oled_colour = 16'b11111_111101_11111; 
		2166: oled_colour = 16'b11111_111111_11111; 
		2167: oled_colour = 16'b10111_111100_11111; 
		2168: oled_colour = 16'b01101_101101_11110; 
		2169: oled_colour = 16'b00111_011101_11001; 
		2170: oled_colour = 16'b00101_010011_10111; 
		2171: oled_colour = 16'b00001_100000_10000; 
		2172: oled_colour = 16'b00001_000001_00001; 
		2173: oled_colour = 16'b00001_000001_00001; 
		2174: oled_colour = 16'b00001_000001_00001; 
		2175: oled_colour = 16'b00001_000001_00001; 
		2176: oled_colour = 16'b00001_000001_00001; 
		2177: oled_colour = 16'b00001_000001_00001; 
		2178: oled_colour = 16'b00001_000001_00001; 
		2179: oled_colour = 16'b00001_000001_00001; 
		2180: oled_colour = 16'b00001_000001_00001; 
		2181: oled_colour = 16'b00001_000001_00001; 
		2182: oled_colour = 16'b00001_000001_00001; 
		2183: oled_colour = 16'b00001_000001_00001; 
		2184: oled_colour = 16'b00001_000001_00001; 
		2185: oled_colour = 16'b00001_000001_00001; 
		2186: oled_colour = 16'b00001_000001_00001; 
		2187: oled_colour = 16'b00001_000001_00001; 
		2188: oled_colour = 16'b00001_000001_00001; 
		2189: oled_colour = 16'b00001_000001_00001; 
		2190: oled_colour = 16'b00001_000001_00001; 
		2191: oled_colour = 16'b00001_000001_00001; 
		2192: oled_colour = 16'b00001_000001_00001; 
		2193: oled_colour = 16'b00001_000001_00001; 
		2194: oled_colour = 16'b00001_000001_00001; 
		2195: oled_colour = 16'b00001_000001_00001; 
		2196: oled_colour = 16'b00001_000001_00001; 
		2197: oled_colour = 16'b00001_000001_00001; 
		2198: oled_colour = 16'b00001_000001_00001; 
		2199: oled_colour = 16'b00001_000001_00001; 
		2200: oled_colour = 16'b00001_000001_00001; 
		2201: oled_colour = 16'b00001_000001_00001; 
		2202: oled_colour = 16'b00001_000001_00001; 
		2203: oled_colour = 16'b00001_000001_00001; 
		2204: oled_colour = 16'b00001_000001_00001; 
		2205: oled_colour = 16'b00001_000001_00001; 
		2206: oled_colour = 16'b00001_000001_00001; 
		2207: oled_colour = 16'b00001_000001_00001; 
		2208: oled_colour = 16'b00001_000001_00001; 
		2209: oled_colour = 16'b00001_000001_00001; 
		2210: oled_colour = 16'b00001_000001_00001; 
		2211: oled_colour = 16'b00001_000001_00001; 
		2212: oled_colour = 16'b00001_000001_00001; 
		2213: oled_colour = 16'b00001_000001_00001; 
		2214: oled_colour = 16'b00001_000001_00001; 
		2215: oled_colour = 16'b00001_000001_00001; 
		2216: oled_colour = 16'b00001_000001_00001; 
		2217: oled_colour = 16'b00001_000001_00001; 
		2218: oled_colour = 16'b00001_000001_00001; 
		2219: oled_colour = 16'b00001_000001_00001; 
		2220: oled_colour = 16'b00001_000001_00001; 
		2221: oled_colour = 16'b00001_000001_00001; 
		2222: oled_colour = 16'b00001_000001_00001; 
		2223: oled_colour = 16'b00001_000001_00001; 
		2224: oled_colour = 16'b00001_000001_00001; 
		2225: oled_colour = 16'b00001_000001_00001; 
		2226: oled_colour = 16'b00001_000001_00001; 
		2227: oled_colour = 16'b00001_000001_00001; 
		2228: oled_colour = 16'b00001_000001_00001; 
		2229: oled_colour = 16'b00001_000001_00001; 
		2230: oled_colour = 16'b00001_000001_00001; 
		2231: oled_colour = 16'b00001_000001_00001; 
		2232: oled_colour = 16'b00001_000001_00001; 
		2233: oled_colour = 16'b00001_000001_00001; 
		2234: oled_colour = 16'b00001_000001_00001; 
		2235: oled_colour = 16'b00001_000001_00001; 
		2236: oled_colour = 16'b00001_000001_00001; 
		2237: oled_colour = 16'b00001_000001_00001; 
		2238: oled_colour = 16'b00001_000001_00001; 
		2239: oled_colour = 16'b00001_000001_00001; 
		2240: oled_colour = 16'b00001_000001_00001; 
		2241: oled_colour = 16'b00001_000001_00001; 
		2242: oled_colour = 16'b00001_000001_00001; 
		2243: oled_colour = 16'b00001_000001_00001; 
		2244: oled_colour = 16'b00001_000001_00001; 
		2245: oled_colour = 16'b00001_000001_00001; 
		2246: oled_colour = 16'b00001_000001_00001; 
		2247: oled_colour = 16'b00001_000001_00001; 
		2248: oled_colour = 16'b00001_000001_00001; 
		2249: oled_colour = 16'b00001_000001_00001; 
		2250: oled_colour = 16'b00001_000001_00001; 
		2251: oled_colour = 16'b00001_000001_00001; 
		2252: oled_colour = 16'b00001_000001_00001; 
		2253: oled_colour = 16'b11111_111111_00001; 
		2254: oled_colour = 16'b00001_000001_11111; 
		2255: oled_colour = 16'b11010_011010_00101; 
		2256: oled_colour = 16'b11101_110111_10000; 
		2257: oled_colour = 16'b11111_111111_11100; 
		2258: oled_colour = 16'b11111_111111_11111; 
		2259: oled_colour = 16'b11111_111111_11111; 
		2260: oled_colour = 16'b11111_111111_11111; 
		2261: oled_colour = 16'b11010_111011_11111; 
		2262: oled_colour = 16'b10010_110001_11101; 
		2263: oled_colour = 16'b01100_101000_11100; 
		2264: oled_colour = 16'b00110_011010_11001; 
		2265: oled_colour = 16'b00001_000001_00001; 
		2266: oled_colour = 16'b00001_000001_00001; 
		2267: oled_colour = 16'b00001_000001_00001; 
		2268: oled_colour = 16'b00001_000001_00001; 
		2269: oled_colour = 16'b00001_000001_00001; 
		2270: oled_colour = 16'b00001_000001_00001; 
		2271: oled_colour = 16'b00001_000001_00001; 
		2272: oled_colour = 16'b00001_000001_00001; 
		2273: oled_colour = 16'b00001_000001_00001; 
		2274: oled_colour = 16'b00001_000001_00001; 
		2275: oled_colour = 16'b00001_000001_00001; 
		2276: oled_colour = 16'b00001_000001_00001; 
		2277: oled_colour = 16'b00001_000001_00001; 
		2278: oled_colour = 16'b00001_000001_00001; 
		2279: oled_colour = 16'b00001_000001_00001; 
		2280: oled_colour = 16'b00001_000001_00001; 
		2281: oled_colour = 16'b00001_000001_00001; 
		2282: oled_colour = 16'b00001_000001_00001; 
		2283: oled_colour = 16'b00001_000001_00001; 
		2284: oled_colour = 16'b00001_000001_00001; 
		2285: oled_colour = 16'b00001_000001_00001; 
		2286: oled_colour = 16'b00001_000001_00001; 
		2287: oled_colour = 16'b00001_000001_00001; 
		2288: oled_colour = 16'b00001_000001_00001; 
		2289: oled_colour = 16'b00001_000001_00001; 
		2290: oled_colour = 16'b00001_000001_00001; 
		2291: oled_colour = 16'b00001_000001_00001; 
		2292: oled_colour = 16'b00001_000001_00001; 
		2293: oled_colour = 16'b00001_000001_00001; 
		2294: oled_colour = 16'b00001_000001_00001; 
		2295: oled_colour = 16'b00001_000001_00001; 
		2296: oled_colour = 16'b00001_000001_00001; 
		2297: oled_colour = 16'b00001_000001_00001; 
		2298: oled_colour = 16'b00001_000001_00001; 
		2299: oled_colour = 16'b00001_000001_00001; 
		2300: oled_colour = 16'b00001_000001_00001; 
		2301: oled_colour = 16'b00001_000001_00001; 
		2302: oled_colour = 16'b00001_000001_00001; 
		2303: oled_colour = 16'b00001_000001_00001; 
		2304: oled_colour = 16'b00001_000001_00001; 
		2305: oled_colour = 16'b00001_000001_00001; 
		2306: oled_colour = 16'b00001_000001_00001; 
		2307: oled_colour = 16'b00001_000001_00001; 
		2308: oled_colour = 16'b00001_000001_00001; 
		2309: oled_colour = 16'b00001_000001_00001; 
		2310: oled_colour = 16'b00001_000001_00001; 
		2311: oled_colour = 16'b00001_000001_00001; 
		2312: oled_colour = 16'b00001_000001_00001; 
		2313: oled_colour = 16'b00001_000001_00001; 
		2314: oled_colour = 16'b00001_000001_00001; 
		2315: oled_colour = 16'b00001_000001_00001; 
		2316: oled_colour = 16'b00001_000001_00001; 
		2317: oled_colour = 16'b00001_000001_00001; 
		2318: oled_colour = 16'b00001_000001_00001; 
		2319: oled_colour = 16'b00001_000001_00001; 
		2320: oled_colour = 16'b00001_000001_00001; 
		2321: oled_colour = 16'b00001_000001_00001; 
		2322: oled_colour = 16'b00001_000001_00001; 
		2323: oled_colour = 16'b00001_000001_00001; 
		2324: oled_colour = 16'b00001_000001_00001; 
		2325: oled_colour = 16'b00001_000001_00001; 
		2326: oled_colour = 16'b00001_000001_00001; 
		2327: oled_colour = 16'b00001_000001_00001; 
		2328: oled_colour = 16'b00001_000001_00001; 
		2329: oled_colour = 16'b00001_000001_00001; 
		2330: oled_colour = 16'b00001_000001_00001; 
		2331: oled_colour = 16'b00001_000001_00001; 
		2332: oled_colour = 16'b00001_000001_00001; 
		2333: oled_colour = 16'b00001_000001_00001; 
		2334: oled_colour = 16'b00001_000001_00001; 
		2335: oled_colour = 16'b00001_000001_00001; 
		2336: oled_colour = 16'b00001_000001_00001; 
		2337: oled_colour = 16'b00001_000001_00001; 
		2338: oled_colour = 16'b00001_000001_00001; 
		2339: oled_colour = 16'b00001_000001_00001; 
		2340: oled_colour = 16'b00001_000001_00001; 
		2341: oled_colour = 16'b00001_000001_00001; 
		2342: oled_colour = 16'b00001_000001_00001; 
		2343: oled_colour = 16'b00001_000001_00001; 
		2344: oled_colour = 16'b00001_000001_00001; 
		2345: oled_colour = 16'b00001_000001_00001; 
		2346: oled_colour = 16'b00001_000001_00001; 
		2347: oled_colour = 16'b00001_000001_00001; 
		2348: oled_colour = 16'b00001_000001_00001; 
		2349: oled_colour = 16'b00001_000001_00001; 
		2350: oled_colour = 16'b00001_000001_00001; 
		2351: oled_colour = 16'b00001_000001_00001; 
		2352: oled_colour = 16'b01110_101001_11101; 
		2353: oled_colour = 16'b10100_110011_11110; 
		2354: oled_colour = 16'b10111_110110_11110; 
		2355: oled_colour = 16'b10110_110100_11101; 
		2356: oled_colour = 16'b10001_101111_11101; 
		2357: oled_colour = 16'b01011_100101_11011; 
		2358: oled_colour = 16'b00001_010011_11000; 
		2359: oled_colour = 16'b00001_000001_00001; 
		2360: oled_colour = 16'b00001_000001_00001; 
		2361: oled_colour = 16'b00001_111111_11111; 
		2362: oled_colour = 16'b00001_000001_00001; 
		2363: oled_colour = 16'b00001_000001_00001; 
		2364: oled_colour = 16'b00001_000001_00001; 
		2365: oled_colour = 16'b00001_000001_00001; 
		2366: oled_colour = 16'b00001_000001_00001; 
		2367: oled_colour = 16'b00001_000001_00001; 
		2368: oled_colour = 16'b00001_000001_00001; 
		2369: oled_colour = 16'b00001_000001_00001; 
		2370: oled_colour = 16'b00001_000001_00001; 
		2371: oled_colour = 16'b00001_000001_00001; 
		2372: oled_colour = 16'b00001_000001_00001; 
		2373: oled_colour = 16'b00001_000001_00001; 
		2374: oled_colour = 16'b00001_000001_00001; 
		2375: oled_colour = 16'b00001_000001_00001; 
		2376: oled_colour = 16'b00001_000001_00001; 
		2377: oled_colour = 16'b00001_000001_00001; 
		2378: oled_colour = 16'b00001_000001_00001; 
		2379: oled_colour = 16'b00001_000001_00001; 
		2380: oled_colour = 16'b00001_000001_00001; 
		2381: oled_colour = 16'b00001_000001_00001; 
		2382: oled_colour = 16'b00001_000001_00001; 
		2383: oled_colour = 16'b00001_000001_00001; 
		2384: oled_colour = 16'b00001_000001_00001; 
		2385: oled_colour = 16'b00001_000001_00001; 
		2386: oled_colour = 16'b00001_000001_00001; 
		2387: oled_colour = 16'b00001_000001_00001; 
		2388: oled_colour = 16'b00001_000001_00001; 
		2389: oled_colour = 16'b00001_000001_00001; 
		2390: oled_colour = 16'b00001_000001_00001; 
		2391: oled_colour = 16'b00001_000001_00001; 
		2392: oled_colour = 16'b00001_000001_00001; 
		2393: oled_colour = 16'b00001_000001_00001; 
		2394: oled_colour = 16'b00001_000001_00001; 
		2395: oled_colour = 16'b00001_000001_00001; 
		2396: oled_colour = 16'b00001_000001_00001; 
		2397: oled_colour = 16'b00001_000001_00001; 
		2398: oled_colour = 16'b00001_000001_00001; 
		2399: oled_colour = 16'b00001_000001_00001; 
		2400: oled_colour = 16'b00001_000001_00001; 
		2401: oled_colour = 16'b00001_000001_00001; 
		2402: oled_colour = 16'b00001_000001_00001; 
		2403: oled_colour = 16'b00001_000001_00001; 
		2404: oled_colour = 16'b00001_000001_00001; 
		2405: oled_colour = 16'b00001_000001_00001; 
		2406: oled_colour = 16'b00001_000001_00001; 
		2407: oled_colour = 16'b00001_000001_00001; 
		2408: oled_colour = 16'b00001_000001_00001; 
		2409: oled_colour = 16'b00001_000001_00001; 
		2410: oled_colour = 16'b00001_000001_00001; 
		2411: oled_colour = 16'b00001_000001_00001; 
		2412: oled_colour = 16'b00001_000001_00001; 
		2413: oled_colour = 16'b00001_000001_00001; 
		2414: oled_colour = 16'b00001_000001_00001; 
		2415: oled_colour = 16'b00001_000001_00001; 
		2416: oled_colour = 16'b00001_000001_00001; 
		2417: oled_colour = 16'b00001_000001_00001; 
		2418: oled_colour = 16'b00001_000001_00001; 
		2419: oled_colour = 16'b00001_000001_00001; 
		2420: oled_colour = 16'b00001_000001_00001; 
		2421: oled_colour = 16'b00001_000001_00001; 
		2422: oled_colour = 16'b00001_000001_00001; 
		2423: oled_colour = 16'b00001_000001_00001; 
		2424: oled_colour = 16'b00001_000001_00001; 
		2425: oled_colour = 16'b00001_000001_00001; 
		2426: oled_colour = 16'b00001_000001_00001; 
		2427: oled_colour = 16'b00001_000001_00001; 
		2428: oled_colour = 16'b00001_000001_00001; 
		2429: oled_colour = 16'b00001_000001_00001; 
		2430: oled_colour = 16'b00001_000001_00001; 
		2431: oled_colour = 16'b00001_000001_00001; 
		2432: oled_colour = 16'b00001_000001_00001; 
		2433: oled_colour = 16'b00001_000001_00001; 
		2434: oled_colour = 16'b00001_000001_00001; 
		2435: oled_colour = 16'b00001_000001_00001; 
		2436: oled_colour = 16'b00001_000001_00001; 
		2437: oled_colour = 16'b00001_000001_00001; 
		2438: oled_colour = 16'b00001_000001_00001; 
		2439: oled_colour = 16'b00001_000001_00001; 
		2440: oled_colour = 16'b00001_000001_00001; 
		2441: oled_colour = 16'b00001_000001_00001; 
		2442: oled_colour = 16'b00001_000001_00001; 
		2443: oled_colour = 16'b00001_000001_00001; 
		2444: oled_colour = 16'b00001_000001_00001; 
		2445: oled_colour = 16'b00001_000001_00001; 
		2446: oled_colour = 16'b00001_000001_00001; 
		2447: oled_colour = 16'b00001_000001_00001; 
		2448: oled_colour = 16'b00001_000001_00001; 
		2449: oled_colour = 16'b00001_000001_00001; 
		2450: oled_colour = 16'b00001_000001_00001; 
		2451: oled_colour = 16'b00001_000001_00001; 
		2452: oled_colour = 16'b00001_000001_00001; 
		2453: oled_colour = 16'b00001_000001_00001; 
		2454: oled_colour = 16'b00001_000001_00001; 
		2455: oled_colour = 16'b11111_111111_11111; 
		2456: oled_colour = 16'b01011_010110_10110; 
		2457: oled_colour = 16'b00001_000001_00001; 
		2458: oled_colour = 16'b00001_000001_00001; 
		2459: oled_colour = 16'b00001_000001_00001; 
		2460: oled_colour = 16'b00001_000001_00001; 
		2461: oled_colour = 16'b00001_000001_00001; 
		2462: oled_colour = 16'b00001_000001_00001; 
		2463: oled_colour = 16'b00001_000001_00001; 
		2464: oled_colour = 16'b00001_000001_00001; 
		2465: oled_colour = 16'b00001_000001_00001; 
		2466: oled_colour = 16'b00001_000001_00001; 
		2467: oled_colour = 16'b00001_000001_00001; 
		2468: oled_colour = 16'b00001_000001_00001; 
		2469: oled_colour = 16'b00001_000001_00001; 
		2470: oled_colour = 16'b00001_000001_00001; 
		2471: oled_colour = 16'b00001_000001_00001; 
		2472: oled_colour = 16'b00001_000001_00001; 
		2473: oled_colour = 16'b00001_000001_00001; 
		2474: oled_colour = 16'b00001_000001_00001; 
		2475: oled_colour = 16'b00001_000001_00001; 
		2476: oled_colour = 16'b00001_000001_00001; 
		2477: oled_colour = 16'b00001_000001_00001; 
		2478: oled_colour = 16'b00001_000001_00001; 
		2479: oled_colour = 16'b00001_000001_00001; 
		2480: oled_colour = 16'b00001_000001_00001; 
		2481: oled_colour = 16'b00001_000001_00001; 
		2482: oled_colour = 16'b00001_000001_00001; 
		2483: oled_colour = 16'b00001_000001_00001; 
		2484: oled_colour = 16'b00001_000001_00001; 
		2485: oled_colour = 16'b00001_000001_00001; 
		2486: oled_colour = 16'b00001_000001_00001; 
		2487: oled_colour = 16'b00001_000001_00001; 
		2488: oled_colour = 16'b00001_000001_00001; 
		2489: oled_colour = 16'b00001_000001_00001; 
		2490: oled_colour = 16'b00001_000001_00001; 
		2491: oled_colour = 16'b00001_000001_00001; 
		2492: oled_colour = 16'b00001_000001_00001; 
		2493: oled_colour = 16'b00001_000001_00001; 
		2494: oled_colour = 16'b00001_000001_00001; 
		2495: oled_colour = 16'b00001_000001_00001; 
		2496: oled_colour = 16'b00001_000001_00001; 
		2497: oled_colour = 16'b00001_000001_00001; 
		2498: oled_colour = 16'b00001_000001_00001; 
		2499: oled_colour = 16'b00001_000001_00001; 
		2500: oled_colour = 16'b00001_000001_00001; 
		2501: oled_colour = 16'b00001_000001_00001; 
		2502: oled_colour = 16'b00001_000001_00001; 
		2503: oled_colour = 16'b00001_000001_00001; 
		2504: oled_colour = 16'b00001_000001_00001; 
		2505: oled_colour = 16'b00001_000001_00001; 
		2506: oled_colour = 16'b00001_000001_00001; 
		2507: oled_colour = 16'b00001_000001_00001; 
		2508: oled_colour = 16'b00001_000001_00001; 
		2509: oled_colour = 16'b00001_000001_00001; 
		2510: oled_colour = 16'b00001_000001_00001; 
		2511: oled_colour = 16'b00001_000001_00001; 
		2512: oled_colour = 16'b00001_000001_00001; 
		2513: oled_colour = 16'b00001_000001_00001; 
		2514: oled_colour = 16'b00001_000001_00001; 
		2515: oled_colour = 16'b00001_000001_00001; 
		2516: oled_colour = 16'b00001_000001_00001; 
		2517: oled_colour = 16'b00001_000001_00001; 
		2518: oled_colour = 16'b00001_000001_00001; 
		2519: oled_colour = 16'b00001_000001_00001; 
		2520: oled_colour = 16'b00001_000001_00001; 
		2521: oled_colour = 16'b00001_000001_00001; 
		2522: oled_colour = 16'b00001_000001_00001; 
		2523: oled_colour = 16'b00001_000001_00001; 
		2524: oled_colour = 16'b00001_000001_00001; 
		2525: oled_colour = 16'b00001_000001_00001; 
		2526: oled_colour = 16'b00001_000001_00001; 
		2527: oled_colour = 16'b00001_000001_00001; 
		2528: oled_colour = 16'b00001_000001_00001; 
		2529: oled_colour = 16'b00001_000001_00001; 
		2530: oled_colour = 16'b00001_000001_00001; 
		2531: oled_colour = 16'b00001_000001_00001; 
		2532: oled_colour = 16'b00001_000001_00001; 
		2533: oled_colour = 16'b00001_000001_00001; 
		2534: oled_colour = 16'b00001_000001_00001; 
		2535: oled_colour = 16'b00001_000001_00001; 
		2536: oled_colour = 16'b00001_000001_00001; 
		2537: oled_colour = 16'b00001_000001_00001; 
		2538: oled_colour = 16'b00001_000001_00001; 
		2539: oled_colour = 16'b00001_000001_00001; 
		2540: oled_colour = 16'b00001_000001_00001; 
		2541: oled_colour = 16'b00001_000001_00001; 
		2542: oled_colour = 16'b00001_000001_00001; 
		2543: oled_colour = 16'b00001_000001_00001; 
		2544: oled_colour = 16'b10000_100000_10000; 
		2545: oled_colour = 16'b11111_111111_11111; 
		2546: oled_colour = 16'b00001_000001_00001; 
		2547: oled_colour = 16'b00001_000001_00001; 
		2548: oled_colour = 16'b11111_111111_11111; 
		2549: oled_colour = 16'b10000_100000_11000; 
		2550: oled_colour = 16'b00001_100000_11111; 
		2551: oled_colour = 16'b00001_000001_00001; 
		2552: oled_colour = 16'b00001_000001_00001; 
		2553: oled_colour = 16'b00001_000001_00001; 
		2554: oled_colour = 16'b00001_000001_00001; 
		2555: oled_colour = 16'b00001_000001_00001; 
		2556: oled_colour = 16'b00001_000001_00001; 
		2557: oled_colour = 16'b00001_000001_00001; 
		2558: oled_colour = 16'b00001_000001_00001; 
		2559: oled_colour = 16'b00001_000001_00001; 
		2560: oled_colour = 16'b00001_000001_00001; 
		2561: oled_colour = 16'b00001_000001_00001; 
		2562: oled_colour = 16'b00001_000001_00001; 
		2563: oled_colour = 16'b00001_000001_00001; 
		2564: oled_colour = 16'b00001_000001_00001; 
		2565: oled_colour = 16'b00001_000001_00001; 
		2566: oled_colour = 16'b00001_000001_00001; 
		2567: oled_colour = 16'b00001_000001_00001; 
		2568: oled_colour = 16'b00001_000001_00001; 
		2569: oled_colour = 16'b00001_000001_00001; 
		2570: oled_colour = 16'b00001_000001_00001; 
		2571: oled_colour = 16'b00001_000001_00001; 
		2572: oled_colour = 16'b00001_000001_00001; 
		2573: oled_colour = 16'b00001_000001_00001; 
		2574: oled_colour = 16'b00001_000001_00001; 
		2575: oled_colour = 16'b00001_000001_00001; 
		2576: oled_colour = 16'b00001_000001_00001; 
		2577: oled_colour = 16'b00001_000001_00001; 
		2578: oled_colour = 16'b00001_000001_00001; 
		2579: oled_colour = 16'b00001_000001_00001; 
		2580: oled_colour = 16'b00001_000001_00001; 
		2581: oled_colour = 16'b00001_000001_00001; 
		2582: oled_colour = 16'b00001_000001_00001; 
		2583: oled_colour = 16'b00001_000001_00001; 
		2584: oled_colour = 16'b00001_000001_00001; 
		2585: oled_colour = 16'b00001_000001_00001; 
		2586: oled_colour = 16'b00001_000001_00001; 
		2587: oled_colour = 16'b00001_000001_00001; 
		2588: oled_colour = 16'b00001_000001_00001; 
		2589: oled_colour = 16'b00001_000001_00001; 
		2590: oled_colour = 16'b00001_000001_00001; 
		2591: oled_colour = 16'b00001_000001_00001; 
		2592: oled_colour = 16'b00001_000001_00001; 
		2593: oled_colour = 16'b00001_000001_00001; 
		2594: oled_colour = 16'b00001_000001_00001; 
		2595: oled_colour = 16'b00001_000001_00001; 
		2596: oled_colour = 16'b00001_000001_00001; 
		2597: oled_colour = 16'b00001_000001_00001; 
		2598: oled_colour = 16'b00001_000001_00001; 
		2599: oled_colour = 16'b00001_000001_00001; 
		2600: oled_colour = 16'b00001_000001_00001; 
		2601: oled_colour = 16'b00001_000001_00001; 
		2602: oled_colour = 16'b00001_000001_00001; 
		2603: oled_colour = 16'b00001_000001_00001; 
		2604: oled_colour = 16'b00001_000001_00001; 
		2605: oled_colour = 16'b00001_000001_00001; 
		2606: oled_colour = 16'b00001_000001_00001; 
		2607: oled_colour = 16'b00001_000001_00001; 
		2608: oled_colour = 16'b00001_000001_00001; 
		2609: oled_colour = 16'b00001_000001_00001; 
		2610: oled_colour = 16'b00001_000001_00001; 
		2611: oled_colour = 16'b00001_000001_00001; 
		2612: oled_colour = 16'b00001_000001_00001; 
		2613: oled_colour = 16'b00001_000001_00001; 
		2614: oled_colour = 16'b00001_000001_00001; 
		2615: oled_colour = 16'b00001_000001_00001; 
		2616: oled_colour = 16'b00001_000001_00001; 
		2617: oled_colour = 16'b00001_000001_00001; 
		2618: oled_colour = 16'b00001_000001_00001; 
		2619: oled_colour = 16'b00001_000001_00001; 
		2620: oled_colour = 16'b00001_000001_00001; 
		2621: oled_colour = 16'b00001_000001_00001; 
		2622: oled_colour = 16'b00001_000001_00001; 
		2623: oled_colour = 16'b00001_000001_00001; 
		2624: oled_colour = 16'b00001_000001_00001; 
		2625: oled_colour = 16'b00001_000001_00001; 
		2626: oled_colour = 16'b00001_000001_00001; 
		2627: oled_colour = 16'b00001_000001_00001; 
		2628: oled_colour = 16'b00001_000001_00001; 
		2629: oled_colour = 16'b00001_000001_00001; 
		2630: oled_colour = 16'b00001_000001_00001; 
		2631: oled_colour = 16'b00001_000001_00001; 
		2632: oled_colour = 16'b00001_000001_00001; 
		2633: oled_colour = 16'b00001_000001_00001; 
		2634: oled_colour = 16'b00001_000001_00001; 
		2635: oled_colour = 16'b00001_000001_00001; 
		2636: oled_colour = 16'b00001_000001_00001; 
		2637: oled_colour = 16'b00001_000001_00001; 
		2638: oled_colour = 16'b00001_000001_00001; 
		2639: oled_colour = 16'b00001_000001_00001; 
		2640: oled_colour = 16'b00001_000001_00001; 
		2641: oled_colour = 16'b00001_000001_00001; 
		2642: oled_colour = 16'b00001_000001_00001; 
		2643: oled_colour = 16'b00001_000001_00001; 
		2644: oled_colour = 16'b00001_000001_00001; 
		2645: oled_colour = 16'b00001_000001_00001; 
		2646: oled_colour = 16'b00001_000001_00001; 
		2647: oled_colour = 16'b00001_000001_00001; 
		2648: oled_colour = 16'b00001_000001_00001; 
		2649: oled_colour = 16'b00001_000001_00001; 
		2650: oled_colour = 16'b00001_000001_00001; 
		2651: oled_colour = 16'b00001_000001_00001; 
		2652: oled_colour = 16'b00001_000001_00001; 
		2653: oled_colour = 16'b00001_000001_00001; 
		2654: oled_colour = 16'b00001_000001_00001; 
		2655: oled_colour = 16'b00001_000001_00001; 
		2656: oled_colour = 16'b00001_000001_00001; 
		2657: oled_colour = 16'b00001_000001_00001; 
		2658: oled_colour = 16'b00001_000001_00001; 
		2659: oled_colour = 16'b00001_000001_00001; 
		2660: oled_colour = 16'b00001_000001_00001; 
		2661: oled_colour = 16'b00001_000001_00001; 
		2662: oled_colour = 16'b00001_000001_00001; 
		2663: oled_colour = 16'b00001_000001_00001; 
		2664: oled_colour = 16'b00001_000001_00001; 
		2665: oled_colour = 16'b00001_000001_00001; 
		2666: oled_colour = 16'b00001_000001_00001; 
		2667: oled_colour = 16'b00001_000001_00001; 
		2668: oled_colour = 16'b00001_000001_00001; 
		2669: oled_colour = 16'b00001_000001_00001; 
		2670: oled_colour = 16'b00001_000001_00001; 
		2671: oled_colour = 16'b00001_000001_00001; 
		2672: oled_colour = 16'b00001_000001_00001; 
		2673: oled_colour = 16'b00001_000001_00001; 
		2674: oled_colour = 16'b00001_000001_00001; 
		2675: oled_colour = 16'b00001_000001_00001; 
		2676: oled_colour = 16'b00001_000001_00001; 
		2677: oled_colour = 16'b00001_000001_00001; 
		2678: oled_colour = 16'b00001_000001_00001; 
		2679: oled_colour = 16'b00001_000001_00001; 
		2680: oled_colour = 16'b00001_000001_00001; 
		2681: oled_colour = 16'b00001_000001_00001; 
		2682: oled_colour = 16'b00001_000001_00001; 
		2683: oled_colour = 16'b00001_000001_00001; 
		2684: oled_colour = 16'b00001_000001_00001; 
		2685: oled_colour = 16'b00001_000001_00001; 
		2686: oled_colour = 16'b00001_000001_00001; 
		2687: oled_colour = 16'b00001_000001_00001; 
		2688: oled_colour = 16'b00001_000001_00001; 
		2689: oled_colour = 16'b00001_000001_00001; 
		2690: oled_colour = 16'b00001_000001_00001; 
		2691: oled_colour = 16'b00001_000001_00001; 
		2692: oled_colour = 16'b00001_000001_00001; 
		2693: oled_colour = 16'b00001_000001_00001; 
		2694: oled_colour = 16'b00001_000001_00001; 
		2695: oled_colour = 16'b00001_000001_00001; 
		2696: oled_colour = 16'b00001_000001_00001; 
		2697: oled_colour = 16'b00001_000001_00001; 
		2698: oled_colour = 16'b00001_000001_00001; 
		2699: oled_colour = 16'b00001_000001_00001; 
		2700: oled_colour = 16'b00001_000001_00001; 
		2701: oled_colour = 16'b00001_000001_00001; 
		2702: oled_colour = 16'b00001_000001_00001; 
		2703: oled_colour = 16'b00001_000001_00001; 
		2704: oled_colour = 16'b00001_000001_00001; 
		2705: oled_colour = 16'b00001_000001_00001; 
		2706: oled_colour = 16'b00001_000001_00001; 
		2707: oled_colour = 16'b00001_000001_00001; 
		2708: oled_colour = 16'b00001_000001_00001; 
		2709: oled_colour = 16'b00001_000001_00001; 
		2710: oled_colour = 16'b00001_000001_00001; 
		2711: oled_colour = 16'b00001_000001_00001; 
		2712: oled_colour = 16'b00001_000001_00001; 
		2713: oled_colour = 16'b00001_000001_00001; 
		2714: oled_colour = 16'b00001_000001_00001; 
		2715: oled_colour = 16'b00001_000001_00001; 
		2716: oled_colour = 16'b00001_000001_00001; 
		2717: oled_colour = 16'b00001_000001_00001; 
		2718: oled_colour = 16'b00001_000001_00001; 
		2719: oled_colour = 16'b00001_000001_00001; 
		2720: oled_colour = 16'b00001_000001_00001; 
		2721: oled_colour = 16'b00001_000001_00001; 
		2722: oled_colour = 16'b00001_000001_00001; 
		2723: oled_colour = 16'b00001_000001_00001; 
		2724: oled_colour = 16'b00001_000001_00001; 
		2725: oled_colour = 16'b00001_000001_00001; 
		2726: oled_colour = 16'b00001_000001_00001; 
		2727: oled_colour = 16'b00001_000001_00001; 
		2728: oled_colour = 16'b00001_000001_00001; 
		2729: oled_colour = 16'b00001_000001_00001; 
		2730: oled_colour = 16'b00001_000001_00001; 
		2731: oled_colour = 16'b00001_000001_00001; 
		2732: oled_colour = 16'b00001_000001_00001; 
		2733: oled_colour = 16'b00001_000001_00001; 
		2734: oled_colour = 16'b00001_000001_00001; 
		2735: oled_colour = 16'b00001_000001_00001; 
		2736: oled_colour = 16'b00001_000001_00001; 
		2737: oled_colour = 16'b00001_000001_00001; 
		2738: oled_colour = 16'b00001_000001_00001; 
		2739: oled_colour = 16'b00001_000001_00001; 
		2740: oled_colour = 16'b00001_000001_00001; 
		2741: oled_colour = 16'b00001_000001_00001; 
		2742: oled_colour = 16'b00001_000001_00001; 
		2743: oled_colour = 16'b00001_000001_00001; 
		2744: oled_colour = 16'b00001_000001_00001; 
		2745: oled_colour = 16'b00001_000001_00001; 
		2746: oled_colour = 16'b00001_000001_00001; 
		2747: oled_colour = 16'b00001_000001_00001; 
		2748: oled_colour = 16'b00001_000001_00001; 
		2749: oled_colour = 16'b00001_000001_00001; 
		2750: oled_colour = 16'b00001_000001_00001; 
		2751: oled_colour = 16'b00001_000001_00001; 
		2752: oled_colour = 16'b00001_000001_00001; 
		2753: oled_colour = 16'b00001_000001_00001; 
		2754: oled_colour = 16'b00001_000001_00001; 
		2755: oled_colour = 16'b00001_000001_00001; 
		2756: oled_colour = 16'b00001_000001_00001; 
		2757: oled_colour = 16'b00001_000001_00001; 
		2758: oled_colour = 16'b00001_000001_00001; 
		2759: oled_colour = 16'b00001_000001_00001; 
		2760: oled_colour = 16'b00001_000001_00001; 
		2761: oled_colour = 16'b00001_000001_00001; 
		2762: oled_colour = 16'b00001_000001_00001; 
		2763: oled_colour = 16'b00001_000001_00001; 
		2764: oled_colour = 16'b00001_000001_00001; 
		2765: oled_colour = 16'b00001_000001_00001; 
		2766: oled_colour = 16'b00001_000001_00001; 
		2767: oled_colour = 16'b00001_000001_00001; 
		2768: oled_colour = 16'b00001_000001_00001; 
		2769: oled_colour = 16'b00001_000001_00001; 
		2770: oled_colour = 16'b00001_000001_00001; 
		2771: oled_colour = 16'b00001_000001_00001; 
		2772: oled_colour = 16'b00001_000001_00001; 
		2773: oled_colour = 16'b00001_000001_00001; 
		2774: oled_colour = 16'b00001_000001_00001; 
		2775: oled_colour = 16'b00001_000001_00001; 
		2776: oled_colour = 16'b00001_000001_00001; 
		2777: oled_colour = 16'b00001_000001_00001; 
		2778: oled_colour = 16'b00001_000001_00001; 
		2779: oled_colour = 16'b00001_000001_00001; 
		2780: oled_colour = 16'b00001_000001_00001; 
		2781: oled_colour = 16'b00001_000001_00001; 
		2782: oled_colour = 16'b00001_000001_00001; 
		2783: oled_colour = 16'b00001_000001_00001; 
		2784: oled_colour = 16'b00001_000001_00001; 
		2785: oled_colour = 16'b00001_000001_00001; 
		2786: oled_colour = 16'b00001_000001_00001; 
		2787: oled_colour = 16'b00001_000001_00001; 
		2788: oled_colour = 16'b00001_000001_00001; 
		2789: oled_colour = 16'b00001_000001_00001; 
		2790: oled_colour = 16'b00001_000001_00001; 
		2791: oled_colour = 16'b00001_000001_00001; 
		2792: oled_colour = 16'b00001_000001_00001; 
		2793: oled_colour = 16'b00001_000001_00001; 
		2794: oled_colour = 16'b00001_000001_00001; 
		2795: oled_colour = 16'b00001_000001_00001; 
		2796: oled_colour = 16'b00001_000001_00001; 
		2797: oled_colour = 16'b00001_000001_00001; 
		2798: oled_colour = 16'b00001_000001_00001; 
		2799: oled_colour = 16'b00001_000001_00001; 
		2800: oled_colour = 16'b00001_000001_00001; 
		2801: oled_colour = 16'b00001_000001_00001; 
		2802: oled_colour = 16'b00001_000001_00001; 
		2803: oled_colour = 16'b00001_000001_00001; 
		2804: oled_colour = 16'b00001_000001_00001; 
		2805: oled_colour = 16'b00001_000001_00001; 
		2806: oled_colour = 16'b00001_000001_00001; 
		2807: oled_colour = 16'b00001_000001_00001; 
		2808: oled_colour = 16'b00001_000001_00001; 
		2809: oled_colour = 16'b00001_000001_00001; 
		2810: oled_colour = 16'b00001_000001_00001; 
		2811: oled_colour = 16'b00001_000001_00001; 
		2812: oled_colour = 16'b00001_000001_00001; 
		2813: oled_colour = 16'b00001_000001_00001; 
		2814: oled_colour = 16'b00001_000001_00001; 
		2815: oled_colour = 16'b00001_000001_00001; 
		2816: oled_colour = 16'b00001_000001_00001; 
		2817: oled_colour = 16'b00001_000001_00001; 
		2818: oled_colour = 16'b00001_000001_00001; 
		2819: oled_colour = 16'b00001_000001_00001; 
		2820: oled_colour = 16'b00001_000001_00001; 
		2821: oled_colour = 16'b00001_000001_00001; 
		2822: oled_colour = 16'b00001_000001_00001; 
		2823: oled_colour = 16'b00001_000001_00001; 
		2824: oled_colour = 16'b00001_000001_00001; 
		2825: oled_colour = 16'b00001_000001_00001; 
		2826: oled_colour = 16'b00001_000001_00001; 
		2827: oled_colour = 16'b00001_000001_00001; 
		2828: oled_colour = 16'b00001_000001_00001; 
		2829: oled_colour = 16'b00001_000001_00001; 
		2830: oled_colour = 16'b00001_000001_00001; 
		2831: oled_colour = 16'b00001_000001_00001; 
		2832: oled_colour = 16'b00001_000001_00001; 
		2833: oled_colour = 16'b00001_000001_00001; 
		2834: oled_colour = 16'b00001_000001_00001; 
		2835: oled_colour = 16'b00001_000001_00001; 
		2836: oled_colour = 16'b00001_000001_00001; 
		2837: oled_colour = 16'b00001_000001_00001; 
		2838: oled_colour = 16'b00001_000001_00001; 
		2839: oled_colour = 16'b00001_000001_00001; 
		2840: oled_colour = 16'b00001_000001_00001; 
		2841: oled_colour = 16'b00001_000001_00001; 
		2842: oled_colour = 16'b00001_000001_00001; 
		2843: oled_colour = 16'b00001_000001_00001; 
		2844: oled_colour = 16'b00001_000001_00001; 
		2845: oled_colour = 16'b00001_000001_00001; 
		2846: oled_colour = 16'b00001_000001_00001; 
		2847: oled_colour = 16'b00001_000001_00001; 
		2848: oled_colour = 16'b00001_000001_00001; 
		2849: oled_colour = 16'b00001_000001_00001; 
		2850: oled_colour = 16'b00001_000001_00001; 
		2851: oled_colour = 16'b00001_000001_00001; 
		2852: oled_colour = 16'b00001_000001_00001; 
		2853: oled_colour = 16'b00001_000001_00001; 
		2854: oled_colour = 16'b00001_000001_00001; 
		2855: oled_colour = 16'b00001_000001_00001; 
		2856: oled_colour = 16'b00001_000001_00001; 
		2857: oled_colour = 16'b00001_000001_00001; 
		2858: oled_colour = 16'b00001_000001_00001; 
		2859: oled_colour = 16'b00001_000001_00001; 
		2860: oled_colour = 16'b00001_000001_00001; 
		2861: oled_colour = 16'b00001_000001_00001; 
		2862: oled_colour = 16'b00001_000001_00001; 
		2863: oled_colour = 16'b00001_000001_00001; 
		2864: oled_colour = 16'b00001_000001_00001; 
		2865: oled_colour = 16'b00001_000001_00001; 
		2866: oled_colour = 16'b00001_000001_00001; 
		2867: oled_colour = 16'b00001_000001_00001; 
		2868: oled_colour = 16'b00001_000001_00001; 
		2869: oled_colour = 16'b00001_000001_00001; 
		2870: oled_colour = 16'b00001_000001_00001; 
		2871: oled_colour = 16'b00001_000001_00001; 
		2872: oled_colour = 16'b00001_000001_00001; 
		2873: oled_colour = 16'b00001_000001_00001; 
		2874: oled_colour = 16'b00001_000001_00001; 
		2875: oled_colour = 16'b00001_000001_00001; 
		2876: oled_colour = 16'b00001_000001_00001; 
		2877: oled_colour = 16'b00001_000001_00001; 
		2878: oled_colour = 16'b00001_000001_00001; 
		2879: oled_colour = 16'b00001_000001_00001; 
		2880: oled_colour = 16'b00001_000001_00001; 
		2881: oled_colour = 16'b00001_000001_00001; 
		2882: oled_colour = 16'b00001_000001_00001; 
		2883: oled_colour = 16'b00001_000001_00001; 
		2884: oled_colour = 16'b00001_000001_00001; 
		2885: oled_colour = 16'b00001_000001_00001; 
		2886: oled_colour = 16'b00001_000001_00001; 
		2887: oled_colour = 16'b00001_000001_00001; 
		2888: oled_colour = 16'b00001_000001_00001; 
		2889: oled_colour = 16'b00001_000001_00001; 
		2890: oled_colour = 16'b00001_000001_00001; 
		2891: oled_colour = 16'b00001_000001_00001; 
		2892: oled_colour = 16'b00001_000001_00001; 
		2893: oled_colour = 16'b00001_000001_00001; 
		2894: oled_colour = 16'b00001_000001_00001; 
		2895: oled_colour = 16'b00001_000001_00001; 
		2896: oled_colour = 16'b00001_000001_00001; 
		2897: oled_colour = 16'b00001_000001_00001; 
		2898: oled_colour = 16'b00001_000001_00001; 
		2899: oled_colour = 16'b00001_000001_00001; 
		2900: oled_colour = 16'b00001_000001_00001; 
		2901: oled_colour = 16'b00001_000001_00001; 
		2902: oled_colour = 16'b00001_000001_00001; 
		2903: oled_colour = 16'b00001_000001_00001; 
		2904: oled_colour = 16'b00001_000001_00001; 
		2905: oled_colour = 16'b00001_000001_00001; 
		2906: oled_colour = 16'b00001_000001_00001; 
		2907: oled_colour = 16'b00001_000001_00001; 
		2908: oled_colour = 16'b00001_000001_00001; 
		2909: oled_colour = 16'b00001_000001_00001; 
		2910: oled_colour = 16'b00001_000001_00001; 
		2911: oled_colour = 16'b00001_000001_00001; 
		2912: oled_colour = 16'b00001_000001_00001; 
		2913: oled_colour = 16'b00001_000001_00001; 
		2914: oled_colour = 16'b00001_000001_00001; 
		2915: oled_colour = 16'b00001_000001_00001; 
		2916: oled_colour = 16'b00001_000001_00001; 
		2917: oled_colour = 16'b00001_000001_00001; 
		2918: oled_colour = 16'b00001_000001_00001; 
		2919: oled_colour = 16'b00001_000001_00001; 
		2920: oled_colour = 16'b00001_000001_00001; 
		2921: oled_colour = 16'b00001_000001_00001; 
		2922: oled_colour = 16'b00001_000001_00001; 
		2923: oled_colour = 16'b00001_000001_00001; 
		2924: oled_colour = 16'b00001_000001_00001; 
		2925: oled_colour = 16'b00001_000001_00001; 
		2926: oled_colour = 16'b00001_000001_00001; 
		2927: oled_colour = 16'b00001_000001_00001; 
		2928: oled_colour = 16'b00001_000001_00001; 
		2929: oled_colour = 16'b00001_000001_00001; 
		2930: oled_colour = 16'b00001_000001_00001; 
		2931: oled_colour = 16'b00001_000001_00001; 
		2932: oled_colour = 16'b00001_000001_00001; 
		2933: oled_colour = 16'b00001_000001_00001; 
		2934: oled_colour = 16'b00001_000001_00001; 
		2935: oled_colour = 16'b00001_000001_00001; 
		2936: oled_colour = 16'b00001_000001_00001; 
		2937: oled_colour = 16'b00001_000001_00001; 
		2938: oled_colour = 16'b00001_000001_00001; 
		2939: oled_colour = 16'b00001_000001_00001; 
		2940: oled_colour = 16'b00001_000001_00001; 
		2941: oled_colour = 16'b00001_000001_00001; 
		2942: oled_colour = 16'b00001_000001_00001; 
		2943: oled_colour = 16'b00001_000001_00001; 
		2944: oled_colour = 16'b00001_000001_00001; 
		2945: oled_colour = 16'b00001_000001_00001; 
		2946: oled_colour = 16'b00001_000001_00001; 
		2947: oled_colour = 16'b00001_000001_00001; 
		2948: oled_colour = 16'b00001_000001_00001; 
		2949: oled_colour = 16'b00001_000001_00001; 
		2950: oled_colour = 16'b00001_000001_00001; 
		2951: oled_colour = 16'b00001_000001_00001; 
		2952: oled_colour = 16'b00001_000001_00001; 
		2953: oled_colour = 16'b00001_000001_00001; 
		2954: oled_colour = 16'b00001_000001_00001; 
		2955: oled_colour = 16'b00001_000001_00001; 
		2956: oled_colour = 16'b00001_000001_00001; 
		2957: oled_colour = 16'b00001_000001_00001; 
		2958: oled_colour = 16'b00001_000001_00001; 
		2959: oled_colour = 16'b00001_000001_00001; 
		2960: oled_colour = 16'b00001_000001_00001; 
		2961: oled_colour = 16'b00001_000001_00001; 
		2962: oled_colour = 16'b00001_000001_00001; 
		2963: oled_colour = 16'b00001_000001_00001; 
		2964: oled_colour = 16'b00001_000001_00001; 
		2965: oled_colour = 16'b00001_000001_00001; 
		2966: oled_colour = 16'b00001_000001_00001; 
		2967: oled_colour = 16'b00001_000001_00001; 
		2968: oled_colour = 16'b00001_000001_00001; 
		2969: oled_colour = 16'b00001_000001_00001; 
		2970: oled_colour = 16'b00001_000001_00001; 
		2971: oled_colour = 16'b00001_000001_00001; 
		2972: oled_colour = 16'b00001_000001_00001; 
		2973: oled_colour = 16'b00001_000001_00001; 
		2974: oled_colour = 16'b00001_000001_00001; 
		2975: oled_colour = 16'b00001_000001_00001; 
		2976: oled_colour = 16'b00001_000001_00001; 
		2977: oled_colour = 16'b00001_000001_00001; 
		2978: oled_colour = 16'b00001_000001_00001; 
		2979: oled_colour = 16'b00001_000001_00001; 
		2980: oled_colour = 16'b00001_000001_00001; 
		2981: oled_colour = 16'b00001_000001_00001; 
		2982: oled_colour = 16'b00001_000001_00001; 
		2983: oled_colour = 16'b00001_000001_00001; 
		2984: oled_colour = 16'b00001_000001_00001; 
		2985: oled_colour = 16'b00001_000001_00001; 
		2986: oled_colour = 16'b00001_000001_00001; 
		2987: oled_colour = 16'b00001_000001_00001; 
		2988: oled_colour = 16'b00001_000001_00001; 
		2989: oled_colour = 16'b00001_000001_00001; 
		2990: oled_colour = 16'b00001_000001_00001; 
		2991: oled_colour = 16'b00001_000001_00001; 
		2992: oled_colour = 16'b00001_000001_00001; 
		2993: oled_colour = 16'b00001_000001_00001; 
		2994: oled_colour = 16'b00001_000001_00001; 
		2995: oled_colour = 16'b00001_000001_00001; 
		2996: oled_colour = 16'b00001_000001_00001; 
		2997: oled_colour = 16'b00001_000001_00001; 
		2998: oled_colour = 16'b00001_000001_00001; 
		2999: oled_colour = 16'b00001_000001_00001; 
		3000: oled_colour = 16'b00001_000001_00001; 
		3001: oled_colour = 16'b00001_000001_00001; 
		3002: oled_colour = 16'b00001_000001_00001; 
		3003: oled_colour = 16'b00001_000001_00001; 
		3004: oled_colour = 16'b00001_000001_00001; 
		3005: oled_colour = 16'b00001_000001_00001; 
		3006: oled_colour = 16'b00001_000001_00001; 
		3007: oled_colour = 16'b00001_000001_00001; 
		3008: oled_colour = 16'b00001_000001_00001; 
		3009: oled_colour = 16'b00001_000001_00001; 
		3010: oled_colour = 16'b00001_000001_00001; 
		3011: oled_colour = 16'b00001_000001_00001; 
		3012: oled_colour = 16'b00001_000001_00001; 
		3013: oled_colour = 16'b00001_000001_00001; 
		3014: oled_colour = 16'b00001_000001_00001; 
		3015: oled_colour = 16'b00001_000001_00001; 
		3016: oled_colour = 16'b00001_000001_00001; 
		3017: oled_colour = 16'b00001_000001_00001; 
		3018: oled_colour = 16'b00001_000001_00001; 
		3019: oled_colour = 16'b00001_000001_00001; 
		3020: oled_colour = 16'b00001_000001_00001; 
		3021: oled_colour = 16'b00001_000001_00001; 
		3022: oled_colour = 16'b00001_000001_00001; 
		3023: oled_colour = 16'b00001_000001_00001; 
		3024: oled_colour = 16'b00001_000001_00001; 
		3025: oled_colour = 16'b00001_000001_00001; 
		3026: oled_colour = 16'b00001_000001_00001; 
		3027: oled_colour = 16'b00001_000001_00001; 
		3028: oled_colour = 16'b00001_000001_00001; 
		3029: oled_colour = 16'b00001_000001_00001; 
		3030: oled_colour = 16'b00001_000001_00001; 
		3031: oled_colour = 16'b00001_000001_00001; 
		3032: oled_colour = 16'b00001_000001_00001; 
		3033: oled_colour = 16'b00001_000001_00001; 
		3034: oled_colour = 16'b00001_000001_00001; 
		3035: oled_colour = 16'b00001_000001_00001; 
		3036: oled_colour = 16'b00001_000001_00001; 
		3037: oled_colour = 16'b00001_000001_00001; 
		3038: oled_colour = 16'b00001_000001_00001; 
		3039: oled_colour = 16'b00001_000001_00001; 
		3040: oled_colour = 16'b00001_000001_00001; 
		3041: oled_colour = 16'b00001_000001_00001; 
		3042: oled_colour = 16'b00001_000001_00001; 
		3043: oled_colour = 16'b00001_000001_00001; 
		3044: oled_colour = 16'b00001_000001_00001; 
		3045: oled_colour = 16'b00001_000001_00001; 
		3046: oled_colour = 16'b00001_000001_00001; 
		3047: oled_colour = 16'b00001_000001_00001; 
		3048: oled_colour = 16'b00001_000001_00001; 
		3049: oled_colour = 16'b00001_000001_00001; 
		3050: oled_colour = 16'b00001_000001_00001; 
		3051: oled_colour = 16'b00001_000001_00001; 
		3052: oled_colour = 16'b00001_000001_00001; 
		3053: oled_colour = 16'b00001_000001_00001; 
		3054: oled_colour = 16'b00001_000001_00001; 
		3055: oled_colour = 16'b00001_000001_00001; 
		3056: oled_colour = 16'b00001_000001_00001; 
		3057: oled_colour = 16'b00001_000001_00001; 
		3058: oled_colour = 16'b00001_000001_00001; 
		3059: oled_colour = 16'b00001_000001_00001; 
		3060: oled_colour = 16'b00001_000001_00001; 
		3061: oled_colour = 16'b00001_000001_00001; 
		3062: oled_colour = 16'b00001_000001_00001; 
		3063: oled_colour = 16'b00001_000001_00001; 
		3064: oled_colour = 16'b00001_000001_00001; 
		3065: oled_colour = 16'b00001_000001_00001; 
		3066: oled_colour = 16'b00001_000001_00001; 
		3067: oled_colour = 16'b00001_000001_00001; 
		3068: oled_colour = 16'b00001_000001_00001; 
		3069: oled_colour = 16'b00001_000001_00001; 
		3070: oled_colour = 16'b00001_000001_00001; 
		3071: oled_colour = 16'b00001_000001_00001; 
		3072: oled_colour = 16'b00001_000001_00001; 
		3073: oled_colour = 16'b00001_000001_00001; 
		3074: oled_colour = 16'b00001_000001_00001; 
		3075: oled_colour = 16'b00001_000001_00001; 
		3076: oled_colour = 16'b00001_000001_00001; 
		3077: oled_colour = 16'b00001_000001_00001; 
		3078: oled_colour = 16'b00001_000001_00001; 
		3079: oled_colour = 16'b00001_000001_00001; 
		3080: oled_colour = 16'b00001_000001_00001; 
		3081: oled_colour = 16'b00001_000001_00001; 
		3082: oled_colour = 16'b00001_000001_00001; 
		3083: oled_colour = 16'b00001_000001_00001; 
		3084: oled_colour = 16'b00001_000001_00001; 
		3085: oled_colour = 16'b00001_000001_00001; 
		3086: oled_colour = 16'b00001_000001_00001; 
		3087: oled_colour = 16'b00001_000001_00001; 
		3088: oled_colour = 16'b00001_000001_00001; 
		3089: oled_colour = 16'b00001_000001_00001; 
		3090: oled_colour = 16'b00001_000001_00001; 
		3091: oled_colour = 16'b00001_000001_00001; 
		3092: oled_colour = 16'b00001_000001_00001; 
		3093: oled_colour = 16'b00001_000001_00001; 
		3094: oled_colour = 16'b00001_000001_00001; 
		3095: oled_colour = 16'b00001_000001_00001; 
		3096: oled_colour = 16'b00001_000001_00001; 
		3097: oled_colour = 16'b00001_000001_00001; 
		3098: oled_colour = 16'b00001_000001_00001; 
		3099: oled_colour = 16'b00001_000001_00001; 
		3100: oled_colour = 16'b00001_000001_00001; 
		3101: oled_colour = 16'b00001_000001_00001; 
		3102: oled_colour = 16'b00001_000001_00001; 
		3103: oled_colour = 16'b00001_000001_00001; 
		3104: oled_colour = 16'b00001_000001_00001; 
		3105: oled_colour = 16'b00001_000001_00001; 
		3106: oled_colour = 16'b00001_000001_00001; 
		3107: oled_colour = 16'b00001_000001_00001; 
		3108: oled_colour = 16'b00001_000001_00001; 
		3109: oled_colour = 16'b00001_000001_00001; 
		3110: oled_colour = 16'b00001_000001_00001; 
		3111: oled_colour = 16'b00001_000001_00001; 
		3112: oled_colour = 16'b00001_000001_00001; 
		3113: oled_colour = 16'b00001_000001_00001; 
		3114: oled_colour = 16'b00001_000001_00001; 
		3115: oled_colour = 16'b00001_000001_00001; 
		3116: oled_colour = 16'b00001_000001_00001; 
		3117: oled_colour = 16'b00001_000001_00001; 
		3118: oled_colour = 16'b00001_000001_00001; 
		3119: oled_colour = 16'b00001_000001_00001; 
		3120: oled_colour = 16'b00001_000001_00001; 
		3121: oled_colour = 16'b00001_000001_00001; 
		3122: oled_colour = 16'b00001_000001_00001; 
		3123: oled_colour = 16'b00001_000001_00001; 
		3124: oled_colour = 16'b00001_000001_00001; 
		3125: oled_colour = 16'b00001_000001_00001; 
		3126: oled_colour = 16'b00001_000001_00001; 
		3127: oled_colour = 16'b00001_000001_00001; 
		3128: oled_colour = 16'b00001_000001_00001; 
		3129: oled_colour = 16'b00001_000001_00001; 
		3130: oled_colour = 16'b00001_000001_00001; 
		3131: oled_colour = 16'b00001_000001_00001; 
		3132: oled_colour = 16'b00001_000001_00001; 
		3133: oled_colour = 16'b00001_000001_00001; 
		3134: oled_colour = 16'b00001_000001_00001; 
		3135: oled_colour = 16'b00001_000001_00001; 
		3136: oled_colour = 16'b00001_000001_00001; 
		3137: oled_colour = 16'b00001_000001_00001; 
		3138: oled_colour = 16'b00001_000001_00001; 
		3139: oled_colour = 16'b00001_000001_00001; 
		3140: oled_colour = 16'b00001_000001_00001; 
		3141: oled_colour = 16'b00001_000001_00001; 
		3142: oled_colour = 16'b00001_000001_00001; 
		3143: oled_colour = 16'b00001_000001_00001; 
		3144: oled_colour = 16'b00001_000001_00001; 
		3145: oled_colour = 16'b00001_000001_00001; 
		3146: oled_colour = 16'b00001_000001_00001; 
		3147: oled_colour = 16'b00001_000001_00001; 
		3148: oled_colour = 16'b00001_000001_00001; 
		3149: oled_colour = 16'b00001_000001_00001; 
		3150: oled_colour = 16'b00001_000001_00001; 
		3151: oled_colour = 16'b00001_000001_00001; 
		3152: oled_colour = 16'b00001_000001_00001; 
		3153: oled_colour = 16'b00001_000001_00001; 
		3154: oled_colour = 16'b00001_000001_00001; 
		3155: oled_colour = 16'b00001_000001_00001; 
		3156: oled_colour = 16'b00001_000001_00001; 
		3157: oled_colour = 16'b00001_000001_00001; 
		3158: oled_colour = 16'b00001_000001_00001; 
		3159: oled_colour = 16'b00001_000001_00001; 
		3160: oled_colour = 16'b00001_000001_00001; 
		3161: oled_colour = 16'b00001_000001_00001; 
		3162: oled_colour = 16'b00001_000001_00001; 
		3163: oled_colour = 16'b00001_000001_00001; 
		3164: oled_colour = 16'b00001_000001_00001; 
		3165: oled_colour = 16'b00001_000001_00001; 
		3166: oled_colour = 16'b00001_000001_00001; 
		3167: oled_colour = 16'b00001_000001_00001; 
		3168: oled_colour = 16'b00001_000001_00001; 
		3169: oled_colour = 16'b00001_000001_00001; 
		3170: oled_colour = 16'b00001_000001_00001; 
		3171: oled_colour = 16'b00001_000001_00001; 
		3172: oled_colour = 16'b00001_000001_00001; 
		3173: oled_colour = 16'b00001_000001_00001; 
		3174: oled_colour = 16'b00001_000001_00001; 
		3175: oled_colour = 16'b00001_000001_00001; 
		3176: oled_colour = 16'b00001_000001_00001; 
		3177: oled_colour = 16'b00001_000001_00001; 
		3178: oled_colour = 16'b00001_000001_00001; 
		3179: oled_colour = 16'b00001_000001_00001; 
		3180: oled_colour = 16'b00001_000001_00001; 
		3181: oled_colour = 16'b00001_000001_00001; 
		3182: oled_colour = 16'b00001_000001_00001; 
		3183: oled_colour = 16'b00001_000001_00001; 
		3184: oled_colour = 16'b00001_000001_00001; 
		3185: oled_colour = 16'b00001_000001_00001; 
		3186: oled_colour = 16'b00001_000001_00001; 
		3187: oled_colour = 16'b00001_000001_00001; 
		3188: oled_colour = 16'b00001_000001_00001; 
		3189: oled_colour = 16'b00001_000001_00001; 
		3190: oled_colour = 16'b00001_000001_00001; 
		3191: oled_colour = 16'b00001_000001_00001; 
		3192: oled_colour = 16'b00001_000001_00001; 
		3193: oled_colour = 16'b00001_000001_00001; 
		3194: oled_colour = 16'b00001_000001_00001; 
		3195: oled_colour = 16'b00001_000001_00001; 
		3196: oled_colour = 16'b00001_000001_00001; 
		3197: oled_colour = 16'b00001_000001_00001; 
		3198: oled_colour = 16'b00001_000001_00001; 
		3199: oled_colour = 16'b00001_000001_00001; 
		3200: oled_colour = 16'b00001_000001_00001; 
		3201: oled_colour = 16'b00001_000001_00001; 
		3202: oled_colour = 16'b00001_000001_00001; 
		3203: oled_colour = 16'b00001_000001_00001; 
		3204: oled_colour = 16'b00001_000001_00001; 
		3205: oled_colour = 16'b00001_000001_00001; 
		3206: oled_colour = 16'b00001_000001_00001; 
		3207: oled_colour = 16'b00001_000001_00001; 
		3208: oled_colour = 16'b00001_000001_00001; 
		3209: oled_colour = 16'b00001_000001_00001; 
		3210: oled_colour = 16'b00001_000001_00001; 
		3211: oled_colour = 16'b00001_000001_00001; 
		3212: oled_colour = 16'b00001_000001_00001; 
		3213: oled_colour = 16'b00001_000001_00001; 
		3214: oled_colour = 16'b00001_000001_00001; 
		3215: oled_colour = 16'b00001_000001_00001; 
		3216: oled_colour = 16'b00001_000001_00001; 
		3217: oled_colour = 16'b00001_000001_00001; 
		3218: oled_colour = 16'b00001_000001_00001; 
		3219: oled_colour = 16'b00001_000001_00001; 
		3220: oled_colour = 16'b00001_000001_00001; 
		3221: oled_colour = 16'b00001_000001_00001; 
		3222: oled_colour = 16'b00001_000001_00001; 
		3223: oled_colour = 16'b00001_000001_00001; 
		3224: oled_colour = 16'b00001_000001_00001; 
		3225: oled_colour = 16'b00001_000001_00001; 
		3226: oled_colour = 16'b00001_000001_00001; 
		3227: oled_colour = 16'b00001_000001_00001; 
		3228: oled_colour = 16'b00001_000001_00001; 
		3229: oled_colour = 16'b00001_000001_00001; 
		3230: oled_colour = 16'b00001_000001_00001; 
		3231: oled_colour = 16'b00001_000001_00001; 
		3232: oled_colour = 16'b00001_000001_00001; 
		3233: oled_colour = 16'b00001_000001_00001; 
		3234: oled_colour = 16'b00001_000001_00001; 
		3235: oled_colour = 16'b00001_000001_00001; 
		3236: oled_colour = 16'b00001_000001_00001; 
		3237: oled_colour = 16'b00001_000001_00001; 
		3238: oled_colour = 16'b00001_000001_00001; 
		3239: oled_colour = 16'b00001_000001_00001; 
		3240: oled_colour = 16'b00001_000001_00001; 
		3241: oled_colour = 16'b00001_000001_00001; 
		3242: oled_colour = 16'b00001_000001_00001; 
		3243: oled_colour = 16'b00001_000001_00001; 
		3244: oled_colour = 16'b00001_000001_00001; 
		3245: oled_colour = 16'b00001_000001_00001; 
		3246: oled_colour = 16'b00001_000001_00001; 
		3247: oled_colour = 16'b00001_000001_00001; 
		3248: oled_colour = 16'b00001_000001_00001; 
		3249: oled_colour = 16'b00001_000001_00001; 
		3250: oled_colour = 16'b00001_000001_00001; 
		3251: oled_colour = 16'b00001_000001_00001; 
		3252: oled_colour = 16'b00001_000001_00001; 
		3253: oled_colour = 16'b00001_000001_00001; 
		3254: oled_colour = 16'b00001_000001_00001; 
		3255: oled_colour = 16'b00001_000001_00001; 
		3256: oled_colour = 16'b00001_000001_00001; 
		3257: oled_colour = 16'b00001_000001_00001; 
		3258: oled_colour = 16'b00001_000001_00001; 
		3259: oled_colour = 16'b00001_000001_00001; 
		3260: oled_colour = 16'b00001_000001_00001; 
		3261: oled_colour = 16'b00001_000001_00001; 
		3262: oled_colour = 16'b00001_000001_00001; 
		3263: oled_colour = 16'b00001_000001_00001; 
		3264: oled_colour = 16'b00001_000001_00001; 
		3265: oled_colour = 16'b00001_000001_00001; 
		3266: oled_colour = 16'b00001_000001_00001; 
		3267: oled_colour = 16'b00001_000001_00001; 
		3268: oled_colour = 16'b00001_000001_00001; 
		3269: oled_colour = 16'b00001_000001_00001; 
		3270: oled_colour = 16'b00001_000001_00001; 
		3271: oled_colour = 16'b00001_000001_00001; 
		3272: oled_colour = 16'b00001_000001_00001; 
		3273: oled_colour = 16'b00001_000001_00001; 
		3274: oled_colour = 16'b00001_000001_00001; 
		3275: oled_colour = 16'b00001_000001_00001; 
		3276: oled_colour = 16'b00001_000001_00001; 
		3277: oled_colour = 16'b00001_000001_00001; 
		3278: oled_colour = 16'b00001_000001_00001; 
		3279: oled_colour = 16'b00001_000001_00001; 
		3280: oled_colour = 16'b00001_000001_00001; 
		3281: oled_colour = 16'b00001_000001_00001; 
		3282: oled_colour = 16'b00001_000001_00001; 
		3283: oled_colour = 16'b00001_000001_00001; 
		3284: oled_colour = 16'b00001_000001_00001; 
		3285: oled_colour = 16'b00001_000001_00001; 
		3286: oled_colour = 16'b00001_000001_00001; 
		3287: oled_colour = 16'b00001_000001_00001; 
		3288: oled_colour = 16'b00001_000001_00001; 
		3289: oled_colour = 16'b00001_000001_00001; 
		3290: oled_colour = 16'b00001_000001_00001; 
		3291: oled_colour = 16'b00001_000001_00001; 
		3292: oled_colour = 16'b00001_000001_00001; 
		3293: oled_colour = 16'b00001_000001_00001; 
		3294: oled_colour = 16'b00001_000001_00001; 
		3295: oled_colour = 16'b00001_000001_00001; 
		3296: oled_colour = 16'b00001_000001_00001; 
		3297: oled_colour = 16'b00001_000001_00001; 
		3298: oled_colour = 16'b00001_000001_00001; 
		3299: oled_colour = 16'b00001_000001_00001; 
		3300: oled_colour = 16'b00001_000001_00001; 
		3301: oled_colour = 16'b00001_000001_00001; 
		3302: oled_colour = 16'b00001_000001_00001; 
		3303: oled_colour = 16'b00001_000001_00001; 
		3304: oled_colour = 16'b00001_000001_00001; 
		3305: oled_colour = 16'b00001_000001_00001; 
		3306: oled_colour = 16'b00001_000001_00001; 
		3307: oled_colour = 16'b00001_000001_00001; 
		3308: oled_colour = 16'b00001_000001_00001; 
		3309: oled_colour = 16'b00001_000001_00001; 
		3310: oled_colour = 16'b00001_000001_00001; 
		3311: oled_colour = 16'b00001_000001_00001; 
		3312: oled_colour = 16'b00001_000001_00001; 
		3313: oled_colour = 16'b00001_000001_00001; 
		3314: oled_colour = 16'b00001_000001_00001; 
		3315: oled_colour = 16'b00001_000001_00001; 
		3316: oled_colour = 16'b00001_000001_00001; 
		3317: oled_colour = 16'b00001_000001_00001; 
		3318: oled_colour = 16'b00001_000001_00001; 
		3319: oled_colour = 16'b00001_000001_00001; 
		3320: oled_colour = 16'b00001_000001_00001; 
		3321: oled_colour = 16'b00001_000001_00001; 
		3322: oled_colour = 16'b00001_000001_00001; 
		3323: oled_colour = 16'b00001_000001_00001; 
		3324: oled_colour = 16'b00001_000001_00001; 
		3325: oled_colour = 16'b00001_000001_00001; 
		3326: oled_colour = 16'b00001_000001_00001; 
		3327: oled_colour = 16'b00001_000001_00001; 
		3328: oled_colour = 16'b00001_000001_00001; 
		3329: oled_colour = 16'b00001_000001_00001; 
		3330: oled_colour = 16'b00001_000001_00001; 
		3331: oled_colour = 16'b00001_000001_00001; 
		3332: oled_colour = 16'b00001_000001_00001; 
		3333: oled_colour = 16'b00001_000001_00001; 
		3334: oled_colour = 16'b00001_000001_00001; 
		3335: oled_colour = 16'b00001_000001_00001; 
		3336: oled_colour = 16'b00001_000001_00001; 
		3337: oled_colour = 16'b00001_000001_00001; 
		3338: oled_colour = 16'b00001_000001_00001; 
		3339: oled_colour = 16'b00001_000001_00001; 
		3340: oled_colour = 16'b00001_000001_00001; 
		3341: oled_colour = 16'b00001_000001_00001; 
		3342: oled_colour = 16'b00001_000001_00001; 
		3343: oled_colour = 16'b00001_000001_00001; 
		3344: oled_colour = 16'b00001_000001_00001; 
		3345: oled_colour = 16'b00001_000001_00001; 
		3346: oled_colour = 16'b00001_000001_00001; 
		3347: oled_colour = 16'b00001_000001_00001; 
		3348: oled_colour = 16'b00001_000001_00001; 
		3349: oled_colour = 16'b00001_000001_00001; 
		3350: oled_colour = 16'b00001_000001_00001; 
		3351: oled_colour = 16'b00001_000001_00001; 
		3352: oled_colour = 16'b00001_000001_00001; 
		3353: oled_colour = 16'b00001_000001_00001; 
		3354: oled_colour = 16'b00001_000001_00001; 
		3355: oled_colour = 16'b00001_000001_00001; 
		3356: oled_colour = 16'b00001_000001_00001; 
		3357: oled_colour = 16'b00001_000001_00001; 
		3358: oled_colour = 16'b00001_000001_00001; 
		3359: oled_colour = 16'b00001_000001_00001; 
		3360: oled_colour = 16'b00001_000001_00001; 
		3361: oled_colour = 16'b00001_000001_00001; 
		3362: oled_colour = 16'b00001_000001_00001; 
		3363: oled_colour = 16'b00001_000001_00001; 
		3364: oled_colour = 16'b00001_000001_00001; 
		3365: oled_colour = 16'b00001_000001_00001; 
		3366: oled_colour = 16'b00001_000001_00001; 
		3367: oled_colour = 16'b00001_000001_00001; 
		3368: oled_colour = 16'b00001_000001_00001; 
		3369: oled_colour = 16'b00001_000001_00001; 
		3370: oled_colour = 16'b00001_000001_00001; 
		3371: oled_colour = 16'b00001_000001_00001; 
		3372: oled_colour = 16'b00001_000001_00001; 
		3373: oled_colour = 16'b00001_000001_00001; 
		3374: oled_colour = 16'b00001_000001_00001; 
		3375: oled_colour = 16'b00001_000001_00001; 
		3376: oled_colour = 16'b00001_000001_00001; 
		3377: oled_colour = 16'b00001_000001_00001; 
		3378: oled_colour = 16'b00001_000001_00001; 
		3379: oled_colour = 16'b00001_000001_00001; 
		3380: oled_colour = 16'b00001_000001_00001; 
		3381: oled_colour = 16'b00001_000001_00001; 
		3382: oled_colour = 16'b00001_000001_00001; 
		3383: oled_colour = 16'b00001_000001_00001; 
		3384: oled_colour = 16'b00001_000001_00001; 
		3385: oled_colour = 16'b00001_000001_00001; 
		3386: oled_colour = 16'b00001_000001_00001; 
		3387: oled_colour = 16'b00001_000001_00001; 
		3388: oled_colour = 16'b00001_000001_00001; 
		3389: oled_colour = 16'b00001_000001_00001; 
		3390: oled_colour = 16'b00001_000001_00001; 
		3391: oled_colour = 16'b00001_000001_00001; 
		3392: oled_colour = 16'b00001_000001_00001; 
		3393: oled_colour = 16'b00001_000001_00001; 
		3394: oled_colour = 16'b00001_000001_00001; 
		3395: oled_colour = 16'b00001_000001_00001; 
		3396: oled_colour = 16'b00001_000001_00001; 
		3397: oled_colour = 16'b00001_000001_00001; 
		3398: oled_colour = 16'b00001_000001_00001; 
		3399: oled_colour = 16'b00001_000001_00001; 
		3400: oled_colour = 16'b00001_000001_00001; 
		3401: oled_colour = 16'b00001_000001_00001; 
		3402: oled_colour = 16'b00001_000001_00001; 
		3403: oled_colour = 16'b00001_000001_00001; 
		3404: oled_colour = 16'b00001_000001_00001; 
		3405: oled_colour = 16'b00001_000001_00001; 
		3406: oled_colour = 16'b00001_000001_00001; 
		3407: oled_colour = 16'b00001_000001_00001; 
		3408: oled_colour = 16'b00001_000001_00001; 
		3409: oled_colour = 16'b00001_000001_00001; 
		3410: oled_colour = 16'b00001_000001_00001; 
		3411: oled_colour = 16'b00001_000001_00001; 
		3412: oled_colour = 16'b00001_000001_00001; 
		3413: oled_colour = 16'b00001_000001_00001; 
		3414: oled_colour = 16'b00001_000001_00001; 
		3415: oled_colour = 16'b00001_000001_00001; 
		3416: oled_colour = 16'b00001_000001_00001; 
		3417: oled_colour = 16'b00001_000001_00001; 
		3418: oled_colour = 16'b00001_000001_00001; 
		3419: oled_colour = 16'b00001_000001_00001; 
		3420: oled_colour = 16'b00001_000001_00001; 
		3421: oled_colour = 16'b00001_000001_00001; 
		3422: oled_colour = 16'b00001_000001_00001; 
		3423: oled_colour = 16'b00001_000001_00001; 
		3424: oled_colour = 16'b00001_000001_00001; 
		3425: oled_colour = 16'b00001_000001_00001; 
		3426: oled_colour = 16'b00001_000001_00001; 
		3427: oled_colour = 16'b00001_000001_00001; 
		3428: oled_colour = 16'b00001_000001_00001; 
		3429: oled_colour = 16'b00001_000001_00001; 
		3430: oled_colour = 16'b00001_000001_00001; 
		3431: oled_colour = 16'b00001_000001_00001; 
		3432: oled_colour = 16'b00001_000001_00001; 
		3433: oled_colour = 16'b00001_000001_00001; 
		3434: oled_colour = 16'b00001_000001_00001; 
		3435: oled_colour = 16'b00001_000001_00001; 
		3436: oled_colour = 16'b00001_000001_00001; 
		3437: oled_colour = 16'b00001_000001_00001; 
		3438: oled_colour = 16'b00001_000001_00001; 
		3439: oled_colour = 16'b00001_000001_00001; 
		3440: oled_colour = 16'b00001_000001_00001; 
		3441: oled_colour = 16'b00001_000001_00001; 
		3442: oled_colour = 16'b00001_000001_00001; 
		3443: oled_colour = 16'b00001_000001_00001; 
		3444: oled_colour = 16'b00001_000001_00001; 
		3445: oled_colour = 16'b00001_000001_00001; 
		3446: oled_colour = 16'b00001_000001_00001; 
		3447: oled_colour = 16'b00001_000001_00001; 
		3448: oled_colour = 16'b00001_000001_00001; 
		3449: oled_colour = 16'b00001_000001_00001; 
		3450: oled_colour = 16'b00001_000001_00001; 
		3451: oled_colour = 16'b00001_000001_00001; 
		3452: oled_colour = 16'b00001_000001_00001; 
		3453: oled_colour = 16'b00001_000001_00001; 
		3454: oled_colour = 16'b00001_000001_00001; 
		3455: oled_colour = 16'b00001_000001_00001; 
		3456: oled_colour = 16'b00001_000001_00001; 
		3457: oled_colour = 16'b00001_000001_00001; 
		3458: oled_colour = 16'b00001_000001_00001; 
		3459: oled_colour = 16'b00001_000001_00001; 
		3460: oled_colour = 16'b00001_000001_00001; 
		3461: oled_colour = 16'b00001_000001_00001; 
		3462: oled_colour = 16'b00001_000001_00001; 
		3463: oled_colour = 16'b00001_000001_00001; 
		3464: oled_colour = 16'b00001_000001_00001; 
		3465: oled_colour = 16'b00001_000001_00001; 
		3466: oled_colour = 16'b00001_000001_00001; 
		3467: oled_colour = 16'b00001_000001_00001; 
		3468: oled_colour = 16'b00001_000001_00001; 
		3469: oled_colour = 16'b00001_000001_00001; 
		3470: oled_colour = 16'b00001_000001_00001; 
		3471: oled_colour = 16'b00001_000001_00001; 
		3472: oled_colour = 16'b00001_000001_00001; 
		3473: oled_colour = 16'b00001_000001_00001; 
		3474: oled_colour = 16'b00001_000001_00001; 
		3475: oled_colour = 16'b00001_000001_00001; 
		3476: oled_colour = 16'b00001_000001_00001; 
		3477: oled_colour = 16'b00001_000001_00001; 
		3478: oled_colour = 16'b00001_000001_00001; 
		3479: oled_colour = 16'b00001_000001_00001; 
		3480: oled_colour = 16'b00001_000001_00001; 
		3481: oled_colour = 16'b00001_000001_00001; 
		3482: oled_colour = 16'b00001_000001_00001; 
		3483: oled_colour = 16'b00001_000001_00001; 
		3484: oled_colour = 16'b00001_000001_00001; 
		3485: oled_colour = 16'b00001_000001_00001; 
		3486: oled_colour = 16'b00001_000001_00001; 
		3487: oled_colour = 16'b00001_000001_00001; 
		3488: oled_colour = 16'b00001_000001_00001; 
		3489: oled_colour = 16'b00001_000001_00001; 
		3490: oled_colour = 16'b00001_000001_00001; 
		3491: oled_colour = 16'b00001_000001_00001; 
		3492: oled_colour = 16'b00001_000001_00001; 
		3493: oled_colour = 16'b00001_000001_00001; 
		3494: oled_colour = 16'b00001_000001_00001; 
		3495: oled_colour = 16'b00001_000001_00001; 
		3496: oled_colour = 16'b00001_000001_00001; 
		3497: oled_colour = 16'b00001_000001_00001; 
		3498: oled_colour = 16'b00001_000001_00001; 
		3499: oled_colour = 16'b00001_000001_00001; 
		3500: oled_colour = 16'b00001_000001_00001; 
		3501: oled_colour = 16'b00001_000001_00001; 
		3502: oled_colour = 16'b00001_000001_00001; 
		3503: oled_colour = 16'b00001_000001_00001; 
		3504: oled_colour = 16'b00001_000001_00001; 
		3505: oled_colour = 16'b00001_000001_00001; 
		3506: oled_colour = 16'b00001_000001_00001; 
		3507: oled_colour = 16'b00001_000001_00001; 
		3508: oled_colour = 16'b00001_000001_00001; 
		3509: oled_colour = 16'b00001_000001_00001; 
		3510: oled_colour = 16'b00001_000001_00001; 
		3511: oled_colour = 16'b00001_000001_00001; 
		3512: oled_colour = 16'b00001_000001_00001; 
		3513: oled_colour = 16'b00001_000001_00001; 
		3514: oled_colour = 16'b00001_000001_00001; 
		3515: oled_colour = 16'b00001_000001_00001; 
		3516: oled_colour = 16'b00001_000001_00001; 
		3517: oled_colour = 16'b00001_000001_00001; 
		3518: oled_colour = 16'b00001_000001_00001; 
		3519: oled_colour = 16'b00001_000001_00001; 
		3520: oled_colour = 16'b00001_000001_00001; 
		3521: oled_colour = 16'b00001_000001_00001; 
		3522: oled_colour = 16'b00001_000001_00001; 
		3523: oled_colour = 16'b00001_000001_00001; 
		3524: oled_colour = 16'b00001_000001_00001; 
		3525: oled_colour = 16'b00001_000001_00001; 
		3526: oled_colour = 16'b00001_000001_00001; 
		3527: oled_colour = 16'b00001_000001_00001; 
		3528: oled_colour = 16'b00001_000001_00001; 
		3529: oled_colour = 16'b00001_000001_00001; 
		3530: oled_colour = 16'b00001_000001_00001; 
		3531: oled_colour = 16'b00001_000001_00001; 
		3532: oled_colour = 16'b00001_000001_00001; 
		3533: oled_colour = 16'b00001_000001_00001; 
		3534: oled_colour = 16'b00001_000001_00001; 
		3535: oled_colour = 16'b00001_000001_00001; 
		3536: oled_colour = 16'b00001_000001_00001; 
		3537: oled_colour = 16'b00001_000001_00001; 
		3538: oled_colour = 16'b00001_000001_00001; 
		3539: oled_colour = 16'b00001_000001_00001; 
		3540: oled_colour = 16'b00001_000001_00001; 
		3541: oled_colour = 16'b00001_000001_00001; 
		3542: oled_colour = 16'b00001_000001_00001; 
		3543: oled_colour = 16'b00001_000001_00001; 
		3544: oled_colour = 16'b00001_000001_00001; 
		3545: oled_colour = 16'b00001_000001_00001; 
		3546: oled_colour = 16'b00001_000001_00001; 
		3547: oled_colour = 16'b00001_000001_00001; 
		3548: oled_colour = 16'b00001_000001_00001; 
		3549: oled_colour = 16'b00001_000001_00001; 
		3550: oled_colour = 16'b00001_000001_00001; 
		3551: oled_colour = 16'b00001_000001_00001; 
		3552: oled_colour = 16'b00001_000001_00001; 
		3553: oled_colour = 16'b00001_000001_00001; 
		3554: oled_colour = 16'b00001_000001_00001; 
		3555: oled_colour = 16'b00001_000001_00001; 
		3556: oled_colour = 16'b00001_000001_00001; 
		3557: oled_colour = 16'b00001_000001_00001; 
		3558: oled_colour = 16'b00001_000001_00001; 
		3559: oled_colour = 16'b00001_000001_00001; 
		3560: oled_colour = 16'b00001_000001_00001; 
		3561: oled_colour = 16'b00001_000001_00001; 
		3562: oled_colour = 16'b00001_000001_00001; 
		3563: oled_colour = 16'b00001_000001_00001; 
		3564: oled_colour = 16'b00001_000001_00001; 
		3565: oled_colour = 16'b00001_000001_00001; 
		3566: oled_colour = 16'b00001_000001_00001; 
		3567: oled_colour = 16'b00001_000001_00001; 
		3568: oled_colour = 16'b00001_000001_00001; 
		3569: oled_colour = 16'b00001_000001_00001; 
		3570: oled_colour = 16'b00001_000001_00001; 
		3571: oled_colour = 16'b00001_000001_00001; 
		3572: oled_colour = 16'b00001_000001_00001; 
		3573: oled_colour = 16'b00001_000001_00001; 
		3574: oled_colour = 16'b00001_000001_00001; 
		3575: oled_colour = 16'b00001_000001_00001; 
		3576: oled_colour = 16'b00001_000001_00001; 
		3577: oled_colour = 16'b00001_000001_00001; 
		3578: oled_colour = 16'b00001_000001_00001; 
		3579: oled_colour = 16'b00001_000001_00001; 
		3580: oled_colour = 16'b00001_000001_00001; 
		3581: oled_colour = 16'b00001_000001_00001; 
		3582: oled_colour = 16'b00001_000001_00001; 
		3583: oled_colour = 16'b00001_000001_00001; 
		3584: oled_colour = 16'b00001_000001_00001; 
		3585: oled_colour = 16'b00001_000001_00001; 
		3586: oled_colour = 16'b00001_000001_00001; 
		3587: oled_colour = 16'b00001_000001_00001; 
		3588: oled_colour = 16'b00001_000001_00001; 
		3589: oled_colour = 16'b00001_000001_00001; 
		3590: oled_colour = 16'b00001_000001_00001; 
		3591: oled_colour = 16'b00001_000001_00001; 
		3592: oled_colour = 16'b00001_000001_00001; 
		3593: oled_colour = 16'b00001_000001_00001; 
		3594: oled_colour = 16'b00001_000001_00001; 
		3595: oled_colour = 16'b00001_000001_00001; 
		3596: oled_colour = 16'b00001_000001_00001; 
		3597: oled_colour = 16'b00001_000001_00001; 
		3598: oled_colour = 16'b00001_000001_00001; 
		3599: oled_colour = 16'b00001_000001_00001; 
		3600: oled_colour = 16'b00001_000001_00001; 
		3601: oled_colour = 16'b00001_000001_00001; 
		3602: oled_colour = 16'b00001_000001_00001; 
		3603: oled_colour = 16'b00001_000001_00001; 
		3604: oled_colour = 16'b00001_000001_00001; 
		3605: oled_colour = 16'b00001_000001_00001; 
		3606: oled_colour = 16'b00001_000001_00001; 
		3607: oled_colour = 16'b00001_000001_00001; 
		3608: oled_colour = 16'b00001_000001_00001; 
		3609: oled_colour = 16'b00001_000001_00001; 
		3610: oled_colour = 16'b00001_000001_00001; 
		3611: oled_colour = 16'b00001_000001_00001; 
		3612: oled_colour = 16'b00001_000001_00001; 
		3613: oled_colour = 16'b00001_000001_00001; 
		3614: oled_colour = 16'b00001_000001_00001; 
		3615: oled_colour = 16'b00001_000001_00001; 
		3616: oled_colour = 16'b00001_000001_00001; 
		3617: oled_colour = 16'b00001_000001_00001; 
		3618: oled_colour = 16'b00001_000001_00001; 
		3619: oled_colour = 16'b00001_000001_00001; 
		3620: oled_colour = 16'b00001_000001_00001; 
		3621: oled_colour = 16'b00001_000001_00001; 
		3622: oled_colour = 16'b00001_000001_00001; 
		3623: oled_colour = 16'b00001_000001_00001; 
		3624: oled_colour = 16'b00001_000001_00001; 
		3625: oled_colour = 16'b00001_000001_00001; 
		3626: oled_colour = 16'b00001_000001_00001; 
		3627: oled_colour = 16'b00001_000001_00001; 
		3628: oled_colour = 16'b00001_000001_00001; 
		3629: oled_colour = 16'b00001_000001_00001; 
		3630: oled_colour = 16'b00001_000001_00001; 
		3631: oled_colour = 16'b00001_000001_00001; 
		3632: oled_colour = 16'b00001_000001_00001; 
		3633: oled_colour = 16'b00001_000001_00001; 
		3634: oled_colour = 16'b00001_000001_00001; 
		3635: oled_colour = 16'b00001_000001_00001; 
		3636: oled_colour = 16'b00001_000001_00001; 
		3637: oled_colour = 16'b00001_000001_00001; 
		3638: oled_colour = 16'b00001_000001_00001; 
		3639: oled_colour = 16'b00001_000001_00001; 
		3640: oled_colour = 16'b00001_000001_00001; 
		3641: oled_colour = 16'b00001_000001_00001; 
		3642: oled_colour = 16'b00001_000001_00001; 
		3643: oled_colour = 16'b00001_000001_00001; 
		3644: oled_colour = 16'b00001_000001_00001; 
		3645: oled_colour = 16'b00001_000001_00001; 
		3646: oled_colour = 16'b00001_000001_00001; 
		3647: oled_colour = 16'b00001_000001_00001; 
		3648: oled_colour = 16'b00001_000001_00001; 
		3649: oled_colour = 16'b00001_000001_00001; 
		3650: oled_colour = 16'b00001_000001_00001; 
		3651: oled_colour = 16'b00001_000001_00001; 
		3652: oled_colour = 16'b00001_000001_00001; 
		3653: oled_colour = 16'b00001_000001_00001; 
		3654: oled_colour = 16'b00001_000001_00001; 
		3655: oled_colour = 16'b00001_000001_00001; 
		3656: oled_colour = 16'b00001_000001_00001; 
		3657: oled_colour = 16'b00001_000001_00001; 
		3658: oled_colour = 16'b00001_000001_00001; 
		3659: oled_colour = 16'b00001_000001_00001; 
		3660: oled_colour = 16'b00001_000001_00001; 
		3661: oled_colour = 16'b00001_000001_00001; 
		3662: oled_colour = 16'b00001_000001_00001; 
		3663: oled_colour = 16'b00001_000001_00001; 
		3664: oled_colour = 16'b00001_000001_00001; 
		3665: oled_colour = 16'b00001_000001_00001; 
		3666: oled_colour = 16'b00001_000001_00001; 
		3667: oled_colour = 16'b00001_000001_00001; 
		3668: oled_colour = 16'b00001_000001_00001; 
		3669: oled_colour = 16'b00001_000001_00001; 
		3670: oled_colour = 16'b00001_000001_00001; 
		3671: oled_colour = 16'b00001_000001_00001; 
		3672: oled_colour = 16'b00001_000001_00001; 
		3673: oled_colour = 16'b00001_000001_00001; 
		3674: oled_colour = 16'b00001_000001_00001; 
		3675: oled_colour = 16'b00001_000001_00001; 
		3676: oled_colour = 16'b00001_000001_00001; 
		3677: oled_colour = 16'b00001_000001_00001; 
		3678: oled_colour = 16'b00001_000001_00001; 
		3679: oled_colour = 16'b00001_000001_00001; 
		3680: oled_colour = 16'b00001_000001_00001; 
		3681: oled_colour = 16'b00001_000001_00001; 
		3682: oled_colour = 16'b00001_000001_00001; 
		3683: oled_colour = 16'b00001_000001_00001; 
		3684: oled_colour = 16'b00001_000001_00001; 
		3685: oled_colour = 16'b00001_000001_00001; 
		3686: oled_colour = 16'b00001_000001_00001; 
		3687: oled_colour = 16'b00001_000001_00001; 
		3688: oled_colour = 16'b00001_000001_00001; 
		3689: oled_colour = 16'b00001_000001_00001; 
		3690: oled_colour = 16'b00001_000001_00001; 
		3691: oled_colour = 16'b00001_000001_00001; 
		3692: oled_colour = 16'b00001_000001_00001; 
		3693: oled_colour = 16'b00001_000001_00001; 
		3694: oled_colour = 16'b00001_000001_00001; 
		3695: oled_colour = 16'b00001_000001_00001; 
		3696: oled_colour = 16'b00001_000001_00001; 
		3697: oled_colour = 16'b00001_000001_00001; 
		3698: oled_colour = 16'b00001_000001_00001; 
		3699: oled_colour = 16'b00001_000001_00001; 
		3700: oled_colour = 16'b00001_000001_00001; 
		3701: oled_colour = 16'b00001_000001_00001; 
		3702: oled_colour = 16'b00001_000001_00001; 
		3703: oled_colour = 16'b00001_000001_00001; 
		3704: oled_colour = 16'b00001_000001_00001; 
		3705: oled_colour = 16'b00001_000001_00001; 
		3706: oled_colour = 16'b00001_000001_00001; 
		3707: oled_colour = 16'b00001_000001_00001; 
		3708: oled_colour = 16'b00001_000001_00001; 
		3709: oled_colour = 16'b00001_000001_00001; 
		3710: oled_colour = 16'b00001_000001_00001; 
		3711: oled_colour = 16'b00001_000001_00001; 
		3712: oled_colour = 16'b00001_000001_00001; 
		3713: oled_colour = 16'b00001_000001_00001; 
		3714: oled_colour = 16'b00001_000001_00001; 
		3715: oled_colour = 16'b00001_000001_00001; 
		3716: oled_colour = 16'b00001_000001_00001; 
		3717: oled_colour = 16'b00001_000001_00001; 
		3718: oled_colour = 16'b00001_000001_00001; 
		3719: oled_colour = 16'b00001_000001_00001; 
		3720: oled_colour = 16'b00001_000001_00001; 
		3721: oled_colour = 16'b00001_000001_00001; 
		3722: oled_colour = 16'b00001_000001_00001; 
		3723: oled_colour = 16'b00001_000001_00001; 
		3724: oled_colour = 16'b00001_000001_00001; 
		3725: oled_colour = 16'b00001_000001_00001; 
		3726: oled_colour = 16'b00001_000001_00001; 
		3727: oled_colour = 16'b00001_000001_00001; 
		3728: oled_colour = 16'b00001_000001_00001; 
		3729: oled_colour = 16'b00001_000001_00001; 
		3730: oled_colour = 16'b00001_000001_00001; 
		3731: oled_colour = 16'b00001_000001_00001; 
		3732: oled_colour = 16'b00001_000001_00001; 
		3733: oled_colour = 16'b00001_000001_00001; 
		3734: oled_colour = 16'b00001_000001_00001; 
		3735: oled_colour = 16'b00001_000001_00001; 
		3736: oled_colour = 16'b00001_000001_00001; 
		3737: oled_colour = 16'b00001_000001_00001; 
		3738: oled_colour = 16'b00001_000001_00001; 
		3739: oled_colour = 16'b00001_000001_00001; 
		3740: oled_colour = 16'b00001_000001_00001; 
		3741: oled_colour = 16'b00001_000001_00001; 
		3742: oled_colour = 16'b00001_000001_00001; 
		3743: oled_colour = 16'b00001_000001_00001; 
		3744: oled_colour = 16'b00001_000001_00001; 
		3745: oled_colour = 16'b00001_000001_00001; 
		3746: oled_colour = 16'b00001_000001_00001; 
		3747: oled_colour = 16'b00001_000001_00001; 
		3748: oled_colour = 16'b00001_000001_00001; 
		3749: oled_colour = 16'b00001_000001_00001; 
		3750: oled_colour = 16'b00001_000001_00001; 
		3751: oled_colour = 16'b00001_000001_00001; 
		3752: oled_colour = 16'b00001_000001_00001; 
		3753: oled_colour = 16'b00001_000001_00001; 
		3754: oled_colour = 16'b00001_000001_00001; 
		3755: oled_colour = 16'b00001_000001_00001; 
		3756: oled_colour = 16'b00001_000001_00001; 
		3757: oled_colour = 16'b00001_000001_00001; 
		3758: oled_colour = 16'b00001_000001_00001; 
		3759: oled_colour = 16'b00001_000001_00001; 
		3760: oled_colour = 16'b00001_000001_00001; 
		3761: oled_colour = 16'b00001_000001_00001; 
		3762: oled_colour = 16'b00001_000001_00001; 
		3763: oled_colour = 16'b00001_000001_00001; 
		3764: oled_colour = 16'b00001_000001_00001; 
		3765: oled_colour = 16'b00001_000001_00001; 
		3766: oled_colour = 16'b00001_000001_00001; 
		3767: oled_colour = 16'b00001_000001_00001; 
		3768: oled_colour = 16'b00001_000001_00001; 
		3769: oled_colour = 16'b00001_000001_00001; 
		3770: oled_colour = 16'b00001_000001_00001; 
		3771: oled_colour = 16'b00001_000001_00001; 
		3772: oled_colour = 16'b00001_000001_00001; 
		3773: oled_colour = 16'b00001_000001_00001; 
		3774: oled_colour = 16'b00001_000001_00001; 
		3775: oled_colour = 16'b00001_000001_00001; 
		3776: oled_colour = 16'b00001_000001_00001; 
		3777: oled_colour = 16'b00001_000001_00001; 
		3778: oled_colour = 16'b00001_000001_00001; 
		3779: oled_colour = 16'b00001_000001_00001; 
		3780: oled_colour = 16'b00001_000001_00001; 
		3781: oled_colour = 16'b00001_000001_00001; 
		3782: oled_colour = 16'b00001_000001_00001; 
		3783: oled_colour = 16'b00001_000001_00001; 
		3784: oled_colour = 16'b00001_000001_00001; 
		3785: oled_colour = 16'b00001_000001_00001; 
		3786: oled_colour = 16'b00001_000001_00001; 
		3787: oled_colour = 16'b00001_000001_00001; 
		3788: oled_colour = 16'b00001_000001_00001; 
		3789: oled_colour = 16'b00001_000001_00001; 
		3790: oled_colour = 16'b00001_000001_00001; 
		3791: oled_colour = 16'b00001_000001_00001; 
		3792: oled_colour = 16'b00001_000001_00001; 
		3793: oled_colour = 16'b00001_000001_00001; 
		3794: oled_colour = 16'b00001_000001_00001; 
		3795: oled_colour = 16'b00001_000001_00001; 
		3796: oled_colour = 16'b00001_000001_00001; 
		3797: oled_colour = 16'b00001_000001_00001; 
		3798: oled_colour = 16'b00001_000001_00001; 
		3799: oled_colour = 16'b00001_000001_00001; 
		3800: oled_colour = 16'b00001_000001_00001; 
		3801: oled_colour = 16'b00001_000001_00001; 
		3802: oled_colour = 16'b00001_000001_00001; 
		3803: oled_colour = 16'b00001_000001_00001; 
		3804: oled_colour = 16'b00001_000001_00001; 
		3805: oled_colour = 16'b00001_000001_00001; 
		3806: oled_colour = 16'b00001_000001_00001; 
		3807: oled_colour = 16'b00001_000001_00001; 
		3808: oled_colour = 16'b00001_000001_00001; 
		3809: oled_colour = 16'b00001_000001_00001; 
		3810: oled_colour = 16'b00001_000001_00001; 
		3811: oled_colour = 16'b00001_000001_00001; 
		3812: oled_colour = 16'b00001_000001_00001; 
		3813: oled_colour = 16'b00001_000001_00001; 
		3814: oled_colour = 16'b00001_000001_00001; 
		3815: oled_colour = 16'b00001_000001_00001; 
		3816: oled_colour = 16'b00001_000001_00001; 
		3817: oled_colour = 16'b00001_000001_00001; 
		3818: oled_colour = 16'b00001_000001_00001; 
		3819: oled_colour = 16'b00001_000001_00001; 
		3820: oled_colour = 16'b00001_000001_00001; 
		3821: oled_colour = 16'b00001_000001_00001; 
		3822: oled_colour = 16'b00001_000001_00001; 
		3823: oled_colour = 16'b00001_000001_00001; 
		3824: oled_colour = 16'b00001_000001_00001; 
		3825: oled_colour = 16'b00001_000001_00001; 
		3826: oled_colour = 16'b00001_000001_00001; 
		3827: oled_colour = 16'b00001_000001_00001; 
		3828: oled_colour = 16'b00001_000001_00001; 
		3829: oled_colour = 16'b00001_000001_00001; 
		3830: oled_colour = 16'b00001_000001_00001; 
		3831: oled_colour = 16'b00001_000001_00001; 
		3832: oled_colour = 16'b00001_000001_00001; 
		3833: oled_colour = 16'b00001_000001_00001; 
		3834: oled_colour = 16'b00001_000001_00001; 
		3835: oled_colour = 16'b00001_000001_00001; 
		3836: oled_colour = 16'b00001_000001_00001; 
		3837: oled_colour = 16'b00001_000001_00001; 
		3838: oled_colour = 16'b00001_000001_00001; 
		3839: oled_colour = 16'b00001_000001_00001; 
		3840: oled_colour = 16'b00001_000001_00001; 
		3841: oled_colour = 16'b00001_000001_00001; 
		3842: oled_colour = 16'b00001_000001_00001; 
		3843: oled_colour = 16'b00001_000001_00001; 
		3844: oled_colour = 16'b00001_000001_00001; 
		3845: oled_colour = 16'b00001_000001_00001; 
		3846: oled_colour = 16'b00001_000001_00001; 
		3847: oled_colour = 16'b00001_000001_00001; 
		3848: oled_colour = 16'b00001_000001_00001; 
		3849: oled_colour = 16'b00001_000001_00001; 
		3850: oled_colour = 16'b00001_000001_00001; 
		3851: oled_colour = 16'b00001_000001_00001; 
		3852: oled_colour = 16'b00001_000001_00001; 
		3853: oled_colour = 16'b00001_000001_00001; 
		3854: oled_colour = 16'b00001_000001_00001; 
		3855: oled_colour = 16'b00001_000001_00001; 
		3856: oled_colour = 16'b00001_000001_00001; 
		3857: oled_colour = 16'b00001_000001_00001; 
		3858: oled_colour = 16'b00001_000001_00001; 
		3859: oled_colour = 16'b00001_000001_00001; 
		3860: oled_colour = 16'b00001_000001_00001; 
		3861: oled_colour = 16'b00001_000001_00001; 
		3862: oled_colour = 16'b00001_000001_00001; 
		3863: oled_colour = 16'b00001_000001_00001; 
		3864: oled_colour = 16'b00001_000001_00001; 
		3865: oled_colour = 16'b00001_000001_00001; 
		3866: oled_colour = 16'b00001_000001_00001; 
		3867: oled_colour = 16'b00001_000001_00001; 
		3868: oled_colour = 16'b00001_000001_00001; 
		3869: oled_colour = 16'b00001_000001_00001; 
		3870: oled_colour = 16'b00001_000001_00001; 
		3871: oled_colour = 16'b00001_000001_00001; 
		3872: oled_colour = 16'b00001_000001_00001; 
		3873: oled_colour = 16'b00001_000001_00001; 
		3874: oled_colour = 16'b00001_000001_00001; 
		3875: oled_colour = 16'b00001_000001_00001; 
		3876: oled_colour = 16'b00001_000001_00001; 
		3877: oled_colour = 16'b00001_000001_00001; 
		3878: oled_colour = 16'b00001_000001_00001; 
		3879: oled_colour = 16'b00001_000001_00001; 
		3880: oled_colour = 16'b00001_000001_00001; 
		3881: oled_colour = 16'b00001_000001_00001; 
		3882: oled_colour = 16'b00001_000001_00001; 
		3883: oled_colour = 16'b00001_000001_00001; 
		3884: oled_colour = 16'b00001_000001_00001; 
		3885: oled_colour = 16'b00001_000001_00001; 
		3886: oled_colour = 16'b00001_000001_00001; 
		3887: oled_colour = 16'b00001_000001_00001; 
		3888: oled_colour = 16'b00001_000001_00001; 
		3889: oled_colour = 16'b00001_000001_00001; 
		3890: oled_colour = 16'b00001_000001_00001; 
		3891: oled_colour = 16'b00001_000001_00001; 
		3892: oled_colour = 16'b00001_000001_00001; 
		3893: oled_colour = 16'b00001_000001_00001; 
		3894: oled_colour = 16'b00001_000001_00001; 
		3895: oled_colour = 16'b00001_000001_00001; 
		3896: oled_colour = 16'b00001_000001_00001; 
		3897: oled_colour = 16'b00001_000001_00001; 
		3898: oled_colour = 16'b00001_000001_00001; 
		3899: oled_colour = 16'b00001_000001_00001; 
		3900: oled_colour = 16'b00001_000001_00001; 
		3901: oled_colour = 16'b00001_000001_00001; 
		3902: oled_colour = 16'b00001_000001_00001; 
		3903: oled_colour = 16'b00001_000001_00001; 
		3904: oled_colour = 16'b00001_000001_00001; 
		3905: oled_colour = 16'b00001_000001_00001; 
		3906: oled_colour = 16'b00001_000001_00001; 
		3907: oled_colour = 16'b00001_000001_00001; 
		3908: oled_colour = 16'b00001_000001_00001; 
		3909: oled_colour = 16'b00001_000001_00001; 
		3910: oled_colour = 16'b00001_000001_00001; 
		3911: oled_colour = 16'b00001_000001_00001; 
		3912: oled_colour = 16'b00001_000001_00001; 
		3913: oled_colour = 16'b00001_000001_00001; 
		3914: oled_colour = 16'b00001_000001_00001; 
		3915: oled_colour = 16'b00001_000001_00001; 
		3916: oled_colour = 16'b00001_000001_00001; 
		3917: oled_colour = 16'b00001_000001_00001; 
		3918: oled_colour = 16'b00001_000001_00001; 
		3919: oled_colour = 16'b00001_000001_00001; 
		3920: oled_colour = 16'b00001_000001_00001; 
		3921: oled_colour = 16'b00001_000001_00001; 
		3922: oled_colour = 16'b00001_000001_00001; 
		3923: oled_colour = 16'b00001_000001_00001; 
		3924: oled_colour = 16'b00001_000001_00001; 
		3925: oled_colour = 16'b00001_000001_00001; 
		3926: oled_colour = 16'b00001_000001_00001; 
		3927: oled_colour = 16'b00001_000001_00001; 
		3928: oled_colour = 16'b00001_000001_00001; 
		3929: oled_colour = 16'b00001_000001_00001; 
		3930: oled_colour = 16'b00001_000001_00001; 
		3931: oled_colour = 16'b00001_000001_00001; 
		3932: oled_colour = 16'b00001_000001_00001; 
		3933: oled_colour = 16'b00001_000001_00001; 
		3934: oled_colour = 16'b00001_000001_00001; 
		3935: oled_colour = 16'b00001_000001_00001; 
		3936: oled_colour = 16'b00001_000001_00001; 
		3937: oled_colour = 16'b00001_000001_00001; 
		3938: oled_colour = 16'b00001_000001_00001; 
		3939: oled_colour = 16'b00001_000001_00001; 
		3940: oled_colour = 16'b00001_000001_00001; 
		3941: oled_colour = 16'b00001_000001_00001; 
		3942: oled_colour = 16'b00001_000001_00001; 
		3943: oled_colour = 16'b00001_000001_00001; 
		3944: oled_colour = 16'b00001_000001_00001; 
		3945: oled_colour = 16'b00001_000001_00001; 
		3946: oled_colour = 16'b00001_000001_00001; 
		3947: oled_colour = 16'b00001_000001_00001; 
		3948: oled_colour = 16'b00001_000001_00001; 
		3949: oled_colour = 16'b00001_000001_00001; 
		3950: oled_colour = 16'b00001_000001_00001; 
		3951: oled_colour = 16'b00001_000001_00001; 
		3952: oled_colour = 16'b00001_000001_00001; 
		3953: oled_colour = 16'b00001_000001_00001; 
		3954: oled_colour = 16'b00001_000001_00001; 
		3955: oled_colour = 16'b00001_000001_00001; 
		3956: oled_colour = 16'b00001_000001_00001; 
		3957: oled_colour = 16'b00001_000001_00001; 
		3958: oled_colour = 16'b00001_000001_00001; 
		3959: oled_colour = 16'b00001_000001_00001; 
		3960: oled_colour = 16'b00001_000001_00001; 
		3961: oled_colour = 16'b00001_000001_00001; 
		3962: oled_colour = 16'b00001_000001_00001; 
		3963: oled_colour = 16'b00001_000001_00001; 
		3964: oled_colour = 16'b00001_000001_00001; 
		3965: oled_colour = 16'b00001_000001_00001; 
		3966: oled_colour = 16'b00001_000001_00001; 
		3967: oled_colour = 16'b00001_000001_00001; 
		3968: oled_colour = 16'b00001_000001_00001; 
		3969: oled_colour = 16'b00001_000001_00001; 
		3970: oled_colour = 16'b00001_000001_00001; 
		3971: oled_colour = 16'b00001_000001_00001; 
		3972: oled_colour = 16'b00001_000001_00001; 
		3973: oled_colour = 16'b00001_000001_00001; 
		3974: oled_colour = 16'b00001_000001_00001; 
		3975: oled_colour = 16'b00001_000001_00001; 
		3976: oled_colour = 16'b00001_000001_00001; 
		3977: oled_colour = 16'b00001_000001_00001; 
		3978: oled_colour = 16'b00001_000001_00001; 
		3979: oled_colour = 16'b00001_000001_00001; 
		3980: oled_colour = 16'b00001_000001_00001; 
		3981: oled_colour = 16'b00001_000001_00001; 
		3982: oled_colour = 16'b00001_000001_00001; 
		3983: oled_colour = 16'b00001_000001_00001; 
		3984: oled_colour = 16'b00001_000001_00001; 
		3985: oled_colour = 16'b00001_000001_00001; 
		3986: oled_colour = 16'b00001_000001_00001; 
		3987: oled_colour = 16'b00001_000001_00001; 
		3988: oled_colour = 16'b00001_000001_00001; 
		3989: oled_colour = 16'b00001_000001_00001; 
		3990: oled_colour = 16'b00001_000001_00001; 
		3991: oled_colour = 16'b00001_000001_00001; 
		3992: oled_colour = 16'b00001_000001_00001; 
		3993: oled_colour = 16'b00001_000001_00001; 
		3994: oled_colour = 16'b00001_000001_00001; 
		3995: oled_colour = 16'b00001_000001_00001; 
		3996: oled_colour = 16'b00001_000001_00001; 
		3997: oled_colour = 16'b00001_000001_00001; 
		3998: oled_colour = 16'b00001_000001_00001; 
		3999: oled_colour = 16'b00001_000001_00001; 
		4000: oled_colour = 16'b00001_000001_00001; 
		4001: oled_colour = 16'b00001_000001_00001; 
		4002: oled_colour = 16'b00001_000001_00001; 
		4003: oled_colour = 16'b00001_000001_00001; 
		4004: oled_colour = 16'b00001_000001_00001; 
		4005: oled_colour = 16'b00001_000001_00001; 
		4006: oled_colour = 16'b00001_000001_00001; 
		4007: oled_colour = 16'b00001_000001_00001; 
		4008: oled_colour = 16'b00001_000001_00001; 
		4009: oled_colour = 16'b00001_000001_00001; 
		4010: oled_colour = 16'b00001_000001_00001; 
		4011: oled_colour = 16'b00001_000001_00001; 
		4012: oled_colour = 16'b00001_000001_00001; 
		4013: oled_colour = 16'b00001_000001_00001; 
		4014: oled_colour = 16'b00001_000001_00001; 
		4015: oled_colour = 16'b00001_000001_00001; 
		4016: oled_colour = 16'b00001_000001_00001; 
		4017: oled_colour = 16'b00001_000001_00001; 
		4018: oled_colour = 16'b00001_000001_00001; 
		4019: oled_colour = 16'b00001_000001_00001; 
		4020: oled_colour = 16'b00001_000001_00001; 
		4021: oled_colour = 16'b00001_000001_00001; 
		4022: oled_colour = 16'b00001_000001_00001; 
		4023: oled_colour = 16'b00001_000001_00001; 
		4024: oled_colour = 16'b00001_000001_00001; 
		4025: oled_colour = 16'b00001_000001_00001; 
		4026: oled_colour = 16'b00001_000001_00001; 
		4027: oled_colour = 16'b00001_000001_00001; 
		4028: oled_colour = 16'b00001_000001_00001; 
		4029: oled_colour = 16'b00001_000001_00001; 
		4030: oled_colour = 16'b00001_000001_00001; 
		4031: oled_colour = 16'b00001_000001_00001; 
		4032: oled_colour = 16'b00001_000001_00001; 
		4033: oled_colour = 16'b00001_000001_00001; 
		4034: oled_colour = 16'b00001_000001_00001; 
		4035: oled_colour = 16'b00001_000001_00001; 
		4036: oled_colour = 16'b00001_000001_00001; 
		4037: oled_colour = 16'b00001_000001_00001; 
		4038: oled_colour = 16'b00001_000001_00001; 
		4039: oled_colour = 16'b00001_000001_00001; 
		4040: oled_colour = 16'b00001_000001_00001; 
		4041: oled_colour = 16'b00001_000001_00001; 
		4042: oled_colour = 16'b00001_000001_00001; 
		4043: oled_colour = 16'b00001_000001_00001; 
		4044: oled_colour = 16'b00001_000001_00001; 
		4045: oled_colour = 16'b00001_000001_00001; 
		4046: oled_colour = 16'b00001_000001_00001; 
		4047: oled_colour = 16'b00001_000001_00001; 
		4048: oled_colour = 16'b00001_000001_00001; 
		4049: oled_colour = 16'b00001_000001_00001; 
		4050: oled_colour = 16'b00001_000001_00001; 
		4051: oled_colour = 16'b00001_000001_00001; 
		4052: oled_colour = 16'b00001_000001_00001; 
		4053: oled_colour = 16'b00001_000001_00001; 
		4054: oled_colour = 16'b00001_000001_00001; 
		4055: oled_colour = 16'b00001_000001_00001; 
		4056: oled_colour = 16'b00001_000001_00001; 
		4057: oled_colour = 16'b00001_000001_00001; 
		4058: oled_colour = 16'b00001_000001_00001; 
		4059: oled_colour = 16'b00001_000001_00001; 
		4060: oled_colour = 16'b00001_000001_00001; 
		4061: oled_colour = 16'b00001_000001_00001; 
		4062: oled_colour = 16'b00001_000001_00001; 
		4063: oled_colour = 16'b00001_000001_00001; 
		4064: oled_colour = 16'b00001_000001_00001; 
		4065: oled_colour = 16'b00001_000001_00001; 
		4066: oled_colour = 16'b00001_000001_00001; 
		4067: oled_colour = 16'b00001_000001_00001; 
		4068: oled_colour = 16'b00001_000001_00001; 
		4069: oled_colour = 16'b00001_000001_00001; 
		4070: oled_colour = 16'b00001_000001_00001; 
		4071: oled_colour = 16'b00001_000001_00001; 
		4072: oled_colour = 16'b00001_000001_00001; 
		4073: oled_colour = 16'b00001_000001_00001; 
		4074: oled_colour = 16'b00001_000001_00001; 
		4075: oled_colour = 16'b00001_000001_00001; 
		4076: oled_colour = 16'b00001_000001_00001; 
		4077: oled_colour = 16'b00001_000001_00001; 
		4078: oled_colour = 16'b00001_000001_00001; 
		4079: oled_colour = 16'b00001_000001_00001; 
		4080: oled_colour = 16'b00001_000001_00001; 
		4081: oled_colour = 16'b00001_000001_00001; 
		4082: oled_colour = 16'b00001_000001_00001; 
		4083: oled_colour = 16'b00001_000001_00001; 
		4084: oled_colour = 16'b00001_000001_00001; 
		4085: oled_colour = 16'b00001_000001_00001; 
		4086: oled_colour = 16'b00001_000001_00001; 
		4087: oled_colour = 16'b00001_000001_00001; 
		4088: oled_colour = 16'b00001_000001_00001; 
		4089: oled_colour = 16'b00001_000001_00001; 
		4090: oled_colour = 16'b00001_000001_00001; 
		4091: oled_colour = 16'b00001_000001_00001; 
		4092: oled_colour = 16'b00001_000001_00001; 
		4093: oled_colour = 16'b00001_000001_00001; 
		4094: oled_colour = 16'b00001_000001_00001; 
		4095: oled_colour = 16'b00001_000001_00001; 
		4096: oled_colour = 16'b00001_000001_00001; 
		4097: oled_colour = 16'b00001_000001_00001; 
		4098: oled_colour = 16'b00001_000001_00001; 
		4099: oled_colour = 16'b00001_000001_00001; 
		4100: oled_colour = 16'b00001_000001_00001; 
		4101: oled_colour = 16'b00001_000001_00001; 
		4102: oled_colour = 16'b00001_000001_00001; 
		4103: oled_colour = 16'b00001_000001_00001; 
		4104: oled_colour = 16'b00001_000001_00001; 
		4105: oled_colour = 16'b00001_000001_00001; 
		4106: oled_colour = 16'b00001_000001_00001; 
		4107: oled_colour = 16'b00001_000001_00001; 
		4108: oled_colour = 16'b00001_000001_00001; 
		4109: oled_colour = 16'b00001_000001_00001; 
		4110: oled_colour = 16'b00001_000001_00001; 
		4111: oled_colour = 16'b00001_000001_00001; 
		4112: oled_colour = 16'b00001_000001_00001; 
		4113: oled_colour = 16'b00001_000001_00001; 
		4114: oled_colour = 16'b00001_000001_00001; 
		4115: oled_colour = 16'b00001_000001_00001; 
		4116: oled_colour = 16'b00001_000001_00001; 
		4117: oled_colour = 16'b00001_000001_00001; 
		4118: oled_colour = 16'b00001_000001_00001; 
		4119: oled_colour = 16'b00001_000001_00001; 
		4120: oled_colour = 16'b00001_000001_00001; 
		4121: oled_colour = 16'b00001_000001_00001; 
		4122: oled_colour = 16'b00001_000001_00001; 
		4123: oled_colour = 16'b00001_000001_00001; 
		4124: oled_colour = 16'b00001_000001_00001; 
		4125: oled_colour = 16'b00001_000001_00001; 
		4126: oled_colour = 16'b00001_000001_00001; 
		4127: oled_colour = 16'b00001_000001_00001; 
		4128: oled_colour = 16'b00001_000001_00001; 
		4129: oled_colour = 16'b00001_000001_00001; 
		4130: oled_colour = 16'b00001_000001_00001; 
		4131: oled_colour = 16'b00001_000001_00001; 
		4132: oled_colour = 16'b00001_000001_00001; 
		4133: oled_colour = 16'b00001_000001_00001; 
		4134: oled_colour = 16'b00001_000001_00001; 
		4135: oled_colour = 16'b00001_000001_00001; 
		4136: oled_colour = 16'b00001_000001_00001; 
		4137: oled_colour = 16'b00001_000001_00001; 
		4138: oled_colour = 16'b00001_000001_00001; 
		4139: oled_colour = 16'b00001_000001_00001; 
		4140: oled_colour = 16'b00001_000001_00001; 
		4141: oled_colour = 16'b00001_000001_00001; 
		4142: oled_colour = 16'b00001_000001_00001; 
		4143: oled_colour = 16'b00001_000001_00001; 
		4144: oled_colour = 16'b00001_000001_00001; 
		4145: oled_colour = 16'b00001_000001_00001; 
		4146: oled_colour = 16'b00001_000001_00001; 
		4147: oled_colour = 16'b00001_000001_00001; 
		4148: oled_colour = 16'b00001_000001_00001; 
		4149: oled_colour = 16'b00001_000001_00001; 
		4150: oled_colour = 16'b00001_000001_00001; 
		4151: oled_colour = 16'b00001_000001_00001; 
		4152: oled_colour = 16'b00001_000001_00001; 
		4153: oled_colour = 16'b00001_000001_00001; 
		4154: oled_colour = 16'b00001_000001_00001; 
		4155: oled_colour = 16'b00001_000001_00001; 
		4156: oled_colour = 16'b00001_000001_00001; 
		4157: oled_colour = 16'b00001_000001_00001; 
		4158: oled_colour = 16'b00001_000001_00001; 
		4159: oled_colour = 16'b00001_000001_00001; 
		4160: oled_colour = 16'b00001_000001_00001; 
		4161: oled_colour = 16'b00001_000001_00001; 
		4162: oled_colour = 16'b00001_000001_00001; 
		4163: oled_colour = 16'b00001_000001_00001; 
		4164: oled_colour = 16'b00001_000001_00001; 
		4165: oled_colour = 16'b00001_000001_00001; 
		4166: oled_colour = 16'b00001_000001_00001; 
		4167: oled_colour = 16'b00001_000001_00001; 
		4168: oled_colour = 16'b00001_000001_00001; 
		4169: oled_colour = 16'b00001_000001_00001; 
		4170: oled_colour = 16'b00001_000001_00001; 
		4171: oled_colour = 16'b00001_000001_00001; 
		4172: oled_colour = 16'b00001_000001_00001; 
		4173: oled_colour = 16'b00001_000001_00001; 
		4174: oled_colour = 16'b00001_000001_00001; 
		4175: oled_colour = 16'b00001_000001_00001; 
		4176: oled_colour = 16'b00001_000001_00001; 
		4177: oled_colour = 16'b00001_000001_00001; 
		4178: oled_colour = 16'b00001_000001_00001; 
		4179: oled_colour = 16'b00001_000001_00001; 
		4180: oled_colour = 16'b00001_000001_00001; 
		4181: oled_colour = 16'b00001_000001_00001; 
		4182: oled_colour = 16'b00001_000001_00001; 
		4183: oled_colour = 16'b00001_000001_00001; 
		4184: oled_colour = 16'b00001_000001_00001; 
		4185: oled_colour = 16'b00001_000001_00001; 
		4186: oled_colour = 16'b00001_000001_00001; 
		4187: oled_colour = 16'b00001_000001_00001; 
		4188: oled_colour = 16'b00001_000001_00001; 
		4189: oled_colour = 16'b00001_000001_00001; 
		4190: oled_colour = 16'b00001_000001_00001; 
		4191: oled_colour = 16'b00001_000001_00001; 
		4192: oled_colour = 16'b00001_000001_00001; 
		4193: oled_colour = 16'b00001_000001_00001; 
		4194: oled_colour = 16'b00001_000001_00001; 
		4195: oled_colour = 16'b00001_000001_00001; 
		4196: oled_colour = 16'b00001_000001_00001; 
		4197: oled_colour = 16'b00001_000001_00001; 
		4198: oled_colour = 16'b00001_000001_00001; 
		4199: oled_colour = 16'b00001_000001_00001; 
		4200: oled_colour = 16'b00001_000001_00001; 
		4201: oled_colour = 16'b00001_000001_00001; 
		4202: oled_colour = 16'b00001_000001_00001; 
		4203: oled_colour = 16'b00001_000001_00001; 
		4204: oled_colour = 16'b00001_000001_00001; 
		4205: oled_colour = 16'b00001_000001_00001; 
		4206: oled_colour = 16'b00001_000001_00001; 
		4207: oled_colour = 16'b00001_000001_00001; 
		4208: oled_colour = 16'b00001_000001_00001; 
		4209: oled_colour = 16'b00001_000001_00001; 
		4210: oled_colour = 16'b00001_000001_00001; 
		4211: oled_colour = 16'b00001_000001_00001; 
		4212: oled_colour = 16'b00001_000001_00001; 
		4213: oled_colour = 16'b00001_000001_00001; 
		4214: oled_colour = 16'b00001_000001_00001; 
		4215: oled_colour = 16'b00001_000001_00001; 
		4216: oled_colour = 16'b00001_000001_00001; 
		4217: oled_colour = 16'b00001_000001_00001; 
		4218: oled_colour = 16'b00001_000001_00001; 
		4219: oled_colour = 16'b00001_000001_00001; 
		4220: oled_colour = 16'b00001_000001_00001; 
		4221: oled_colour = 16'b00001_000001_00001; 
		4222: oled_colour = 16'b00001_000001_00001; 
		4223: oled_colour = 16'b00001_000001_00001; 
		4224: oled_colour = 16'b00001_000001_00001; 
		4225: oled_colour = 16'b00001_000001_00001; 
		4226: oled_colour = 16'b00001_000001_00001; 
		4227: oled_colour = 16'b00001_000001_00001; 
		4228: oled_colour = 16'b00001_000001_00001; 
		4229: oled_colour = 16'b00001_000001_00001; 
		4230: oled_colour = 16'b00001_000001_00001; 
		4231: oled_colour = 16'b00001_000001_00001; 
		4232: oled_colour = 16'b00001_000001_00001; 
		4233: oled_colour = 16'b00001_000001_00001; 
		4234: oled_colour = 16'b00001_000001_00001; 
		4235: oled_colour = 16'b00001_000001_00001; 
		4236: oled_colour = 16'b00001_000001_00001; 
		4237: oled_colour = 16'b00001_000001_00001; 
		4238: oled_colour = 16'b00001_000001_00001; 
		4239: oled_colour = 16'b00001_000001_00001; 
		4240: oled_colour = 16'b00001_000001_00001; 
		4241: oled_colour = 16'b00001_000001_00001; 
		4242: oled_colour = 16'b00001_000001_00001; 
		4243: oled_colour = 16'b00001_000001_00001; 
		4244: oled_colour = 16'b00001_000001_00001; 
		4245: oled_colour = 16'b00001_000001_00001; 
		4246: oled_colour = 16'b00001_000001_00001; 
		4247: oled_colour = 16'b00001_000001_00001; 
		4248: oled_colour = 16'b00001_000001_00001; 
		4249: oled_colour = 16'b00001_000001_00001; 
		4250: oled_colour = 16'b00001_000001_00001; 
		4251: oled_colour = 16'b00001_000001_00001; 
		4252: oled_colour = 16'b00001_000001_00001; 
		4253: oled_colour = 16'b00001_000001_00001; 
		4254: oled_colour = 16'b00001_000001_00001; 
		4255: oled_colour = 16'b00001_000001_00001; 
		4256: oled_colour = 16'b00001_000001_00001; 
		4257: oled_colour = 16'b00001_000001_00001; 
		4258: oled_colour = 16'b00001_000001_00001; 
		4259: oled_colour = 16'b00001_000001_00001; 
		4260: oled_colour = 16'b00001_000001_00001; 
		4261: oled_colour = 16'b00001_000001_00001; 
		4262: oled_colour = 16'b00001_000001_00001; 
		4263: oled_colour = 16'b00001_000001_00001; 
		4264: oled_colour = 16'b00001_000001_00001; 
		4265: oled_colour = 16'b00001_000001_00001; 
		4266: oled_colour = 16'b00001_000001_00001; 
		4267: oled_colour = 16'b00001_000001_00001; 
		4268: oled_colour = 16'b00001_000001_00001; 
		4269: oled_colour = 16'b00001_000001_00001; 
		4270: oled_colour = 16'b00001_000001_00001; 
		4271: oled_colour = 16'b00001_000001_00001; 
		4272: oled_colour = 16'b00001_000001_00001; 
		4273: oled_colour = 16'b00001_000001_00001; 
		4274: oled_colour = 16'b00001_000001_00001; 
		4275: oled_colour = 16'b00001_000001_00001; 
		4276: oled_colour = 16'b00001_000001_00001; 
		4277: oled_colour = 16'b00001_000001_00001; 
		4278: oled_colour = 16'b00001_000001_00001; 
		4279: oled_colour = 16'b00001_000001_00001; 
		4280: oled_colour = 16'b00001_000001_00001; 
		4281: oled_colour = 16'b00001_000001_00001; 
		4282: oled_colour = 16'b00001_000001_00001; 
		4283: oled_colour = 16'b00001_000001_00001; 
		4284: oled_colour = 16'b00001_000001_00001; 
		4285: oled_colour = 16'b00001_000001_00001; 
		4286: oled_colour = 16'b00001_000001_00001; 
		4287: oled_colour = 16'b00001_000001_00001; 
		4288: oled_colour = 16'b00001_000001_00001; 
		4289: oled_colour = 16'b00001_000001_00001; 
		4290: oled_colour = 16'b00001_000001_00001; 
		4291: oled_colour = 16'b00001_000001_00001; 
		4292: oled_colour = 16'b00001_000001_00001; 
		4293: oled_colour = 16'b00001_000001_00001; 
		4294: oled_colour = 16'b00001_000001_00001; 
		4295: oled_colour = 16'b00001_000001_00001; 
		4296: oled_colour = 16'b00001_000001_00001; 
		4297: oled_colour = 16'b00001_000001_00001; 
		4298: oled_colour = 16'b00001_000001_00001; 
		4299: oled_colour = 16'b00001_000001_00001; 
		4300: oled_colour = 16'b00001_000001_00001; 
		4301: oled_colour = 16'b00001_000001_00001; 
		4302: oled_colour = 16'b00001_000001_00001; 
		4303: oled_colour = 16'b00001_000001_00001; 
		4304: oled_colour = 16'b00001_000001_00001; 
		4305: oled_colour = 16'b00001_000001_00001; 
		4306: oled_colour = 16'b00001_000001_00001; 
		4307: oled_colour = 16'b00001_000001_00001; 
		4308: oled_colour = 16'b00001_000001_00001; 
		4309: oled_colour = 16'b00001_000001_00001; 
		4310: oled_colour = 16'b00001_000001_00001; 
		4311: oled_colour = 16'b00001_000001_00001; 
		4312: oled_colour = 16'b00001_000001_00001; 
		4313: oled_colour = 16'b00001_000001_00001; 
		4314: oled_colour = 16'b00001_000001_00001; 
		4315: oled_colour = 16'b00001_000001_00001; 
		4316: oled_colour = 16'b00001_000001_00001; 
		4317: oled_colour = 16'b00001_000001_00001; 
		4318: oled_colour = 16'b00001_000001_00001; 
		4319: oled_colour = 16'b00001_000001_00001; 
		4320: oled_colour = 16'b00001_000001_00001; 
		4321: oled_colour = 16'b00001_000001_00001; 
		4322: oled_colour = 16'b00001_000001_00001; 
		4323: oled_colour = 16'b00001_000001_00001; 
		4324: oled_colour = 16'b00001_000001_00001; 
		4325: oled_colour = 16'b00001_000001_00001; 
		4326: oled_colour = 16'b00001_000001_00001; 
		4327: oled_colour = 16'b00001_000001_00001; 
		4328: oled_colour = 16'b00001_000001_00001; 
		4329: oled_colour = 16'b00001_000001_00001; 
		4330: oled_colour = 16'b00001_000001_00001; 
		4331: oled_colour = 16'b00001_000001_00001; 
		4332: oled_colour = 16'b00001_000001_00001; 
		4333: oled_colour = 16'b00001_000001_00001; 
		4334: oled_colour = 16'b00001_000001_00001; 
		4335: oled_colour = 16'b00001_000001_00001; 
		4336: oled_colour = 16'b00001_000001_00001; 
		4337: oled_colour = 16'b00001_000001_00001; 
		4338: oled_colour = 16'b00001_000001_00001; 
		4339: oled_colour = 16'b00001_000001_00001; 
		4340: oled_colour = 16'b00001_000001_00001; 
		4341: oled_colour = 16'b00001_000001_00001; 
		4342: oled_colour = 16'b00001_000001_00001; 
		4343: oled_colour = 16'b00001_000001_00001; 
		4344: oled_colour = 16'b00001_000001_00001; 
		4345: oled_colour = 16'b00001_000001_00001; 
		4346: oled_colour = 16'b00001_000001_00001; 
		4347: oled_colour = 16'b00001_000001_00001; 
		4348: oled_colour = 16'b00001_000001_00001; 
		4349: oled_colour = 16'b00001_000001_00001; 
		4350: oled_colour = 16'b00001_000001_00001; 
		4351: oled_colour = 16'b00001_000001_00001; 
		4352: oled_colour = 16'b00001_000001_00001; 
		4353: oled_colour = 16'b00001_000001_00001; 
		4354: oled_colour = 16'b00001_000001_00001; 
		4355: oled_colour = 16'b00001_000001_00001; 
		4356: oled_colour = 16'b00001_000001_00001; 
		4357: oled_colour = 16'b00001_000001_00001; 
		4358: oled_colour = 16'b00001_000001_00001; 
		4359: oled_colour = 16'b00001_000001_00001; 
		4360: oled_colour = 16'b00001_000001_00001; 
		4361: oled_colour = 16'b00001_000001_00001; 
		4362: oled_colour = 16'b00001_000001_00001; 
		4363: oled_colour = 16'b00001_000001_00001; 
		4364: oled_colour = 16'b00001_000001_00001; 
		4365: oled_colour = 16'b00001_000001_00001; 
		4366: oled_colour = 16'b00001_000001_00001; 
		4367: oled_colour = 16'b00001_000001_00001; 
		4368: oled_colour = 16'b00001_000001_00001; 
		4369: oled_colour = 16'b00001_000001_00001; 
		4370: oled_colour = 16'b00001_000001_00001; 
		4371: oled_colour = 16'b00001_000001_00001; 
		4372: oled_colour = 16'b00001_000001_00001; 
		4373: oled_colour = 16'b00001_000001_00001; 
		4374: oled_colour = 16'b00001_000001_00001; 
		4375: oled_colour = 16'b00001_000001_00001; 
		4376: oled_colour = 16'b00001_000001_00001; 
		4377: oled_colour = 16'b00001_000001_00001; 
		4378: oled_colour = 16'b00001_000001_00001; 
		4379: oled_colour = 16'b00001_000001_00001; 
		4380: oled_colour = 16'b00001_000001_00001; 
		4381: oled_colour = 16'b00001_000001_00001; 
		4382: oled_colour = 16'b00001_000001_00001; 
		4383: oled_colour = 16'b00001_000001_00001; 
		4384: oled_colour = 16'b00001_000001_00001; 
		4385: oled_colour = 16'b00001_000001_00001; 
		4386: oled_colour = 16'b00001_000001_00001; 
		4387: oled_colour = 16'b00001_000001_00001; 
		4388: oled_colour = 16'b00001_000001_00001; 
		4389: oled_colour = 16'b00001_000001_00001; 
		4390: oled_colour = 16'b00001_000001_00001; 
		4391: oled_colour = 16'b00001_000001_00001; 
		4392: oled_colour = 16'b00001_000001_00001; 
		4393: oled_colour = 16'b00001_000001_00001; 
		4394: oled_colour = 16'b00001_000001_00001; 
		4395: oled_colour = 16'b00001_000001_00001; 
		4396: oled_colour = 16'b00001_000001_00001; 
		4397: oled_colour = 16'b00001_000001_00001; 
		4398: oled_colour = 16'b00001_000001_00001; 
		4399: oled_colour = 16'b00001_000001_00001; 
		4400: oled_colour = 16'b00001_000001_00001; 
		4401: oled_colour = 16'b00001_000001_00001; 
		4402: oled_colour = 16'b00001_000001_00001; 
		4403: oled_colour = 16'b00001_000001_00001; 
		4404: oled_colour = 16'b00001_000001_00001; 
		4405: oled_colour = 16'b00001_000001_00001; 
		4406: oled_colour = 16'b00001_000001_00001; 
		4407: oled_colour = 16'b00001_000001_00001; 
		4408: oled_colour = 16'b00001_000001_00001; 
		4409: oled_colour = 16'b00001_000001_00001; 
		4410: oled_colour = 16'b00001_000001_00001; 
		4411: oled_colour = 16'b00001_000001_00001; 
		4412: oled_colour = 16'b00001_000001_00001; 
		4413: oled_colour = 16'b00001_000001_00001; 
		4414: oled_colour = 16'b00001_000001_00001; 
		4415: oled_colour = 16'b00001_000001_00001; 
		4416: oled_colour = 16'b00001_000001_00001; 
		4417: oled_colour = 16'b00001_000001_00001; 
		4418: oled_colour = 16'b00001_000001_00001; 
		4419: oled_colour = 16'b00001_000001_00001; 
		4420: oled_colour = 16'b00001_000001_00001; 
		4421: oled_colour = 16'b00001_000001_00001; 
		4422: oled_colour = 16'b00001_000001_00001; 
		4423: oled_colour = 16'b00001_000001_00001; 
		4424: oled_colour = 16'b00001_000001_00001; 
		4425: oled_colour = 16'b00001_000001_00001; 
		4426: oled_colour = 16'b00001_000001_00001; 
		4427: oled_colour = 16'b00001_000001_00001; 
		4428: oled_colour = 16'b00001_000001_00001; 
		4429: oled_colour = 16'b00001_000001_00001; 
		4430: oled_colour = 16'b00001_000001_00001; 
		4431: oled_colour = 16'b00001_000001_00001; 
		4432: oled_colour = 16'b00001_000001_00001; 
		4433: oled_colour = 16'b00001_000001_00001; 
		4434: oled_colour = 16'b00001_000001_00001; 
		4435: oled_colour = 16'b00001_000001_00001; 
		4436: oled_colour = 16'b00001_000001_00001; 
		4437: oled_colour = 16'b00001_000001_00001; 
		4438: oled_colour = 16'b00001_000001_00001; 
		4439: oled_colour = 16'b00001_000001_00001; 
		4440: oled_colour = 16'b00001_000001_00001; 
		4441: oled_colour = 16'b00001_000001_00001; 
		4442: oled_colour = 16'b00001_000001_00001; 
		4443: oled_colour = 16'b00001_000001_00001; 
		4444: oled_colour = 16'b00001_000001_00001; 
		4445: oled_colour = 16'b00001_000001_00001; 
		4446: oled_colour = 16'b00001_000001_00001; 
		4447: oled_colour = 16'b00001_000001_00001; 
		4448: oled_colour = 16'b00001_000001_00001; 
		4449: oled_colour = 16'b00001_000001_00001; 
		4450: oled_colour = 16'b00001_000001_00001; 
		4451: oled_colour = 16'b00001_000001_00001; 
		4452: oled_colour = 16'b00001_000001_00001; 
		4453: oled_colour = 16'b00001_000001_00001; 
		4454: oled_colour = 16'b00001_000001_00001; 
		4455: oled_colour = 16'b00001_000001_00001; 
		4456: oled_colour = 16'b00001_000001_00001; 
		4457: oled_colour = 16'b00001_000001_00001; 
		4458: oled_colour = 16'b00001_000001_00001; 
		4459: oled_colour = 16'b00001_000001_00001; 
		4460: oled_colour = 16'b00001_000001_00001; 
		4461: oled_colour = 16'b00001_000001_00001; 
		4462: oled_colour = 16'b00001_000001_00001; 
		4463: oled_colour = 16'b00001_000001_00001; 
		4464: oled_colour = 16'b00001_000001_00001; 
		4465: oled_colour = 16'b00001_000001_00001; 
		4466: oled_colour = 16'b00001_000001_00001; 
		4467: oled_colour = 16'b00001_000001_00001; 
		4468: oled_colour = 16'b00001_000001_00001; 
		4469: oled_colour = 16'b00001_000001_00001; 
		4470: oled_colour = 16'b00001_000001_00001; 
		4471: oled_colour = 16'b00001_000001_00001; 
		4472: oled_colour = 16'b00001_000001_00001; 
		4473: oled_colour = 16'b00001_000001_00001; 
		4474: oled_colour = 16'b00001_000001_00001; 
		4475: oled_colour = 16'b00001_000001_00001; 
		4476: oled_colour = 16'b00001_000001_00001; 
		4477: oled_colour = 16'b00001_000001_00001; 
		4478: oled_colour = 16'b00001_000001_00001; 
		4479: oled_colour = 16'b00001_000001_00001; 
		4480: oled_colour = 16'b00001_000001_00001; 
		4481: oled_colour = 16'b00001_000001_00001; 
		4482: oled_colour = 16'b00001_000001_00001; 
		4483: oled_colour = 16'b00001_000001_00001; 
		4484: oled_colour = 16'b00001_000001_00001; 
		4485: oled_colour = 16'b00001_000001_00001; 
		4486: oled_colour = 16'b00001_000001_00001; 
		4487: oled_colour = 16'b00001_000001_00001; 
		4488: oled_colour = 16'b00001_000001_00001; 
		4489: oled_colour = 16'b00001_000001_00001; 
		4490: oled_colour = 16'b00001_000001_00001; 
		4491: oled_colour = 16'b00001_000001_00001; 
		4492: oled_colour = 16'b00001_000001_00001; 
		4493: oled_colour = 16'b00001_000001_00001; 
		4494: oled_colour = 16'b00001_000001_00001; 
		4495: oled_colour = 16'b00001_000001_00001; 
		4496: oled_colour = 16'b00001_000001_00001; 
		4497: oled_colour = 16'b00001_000001_00001; 
		4498: oled_colour = 16'b00001_000001_00001; 
		4499: oled_colour = 16'b00001_000001_00001; 
		4500: oled_colour = 16'b00001_000001_00001; 
		4501: oled_colour = 16'b00001_000001_00001; 
		4502: oled_colour = 16'b00001_000001_00001; 
		4503: oled_colour = 16'b00001_000001_00001; 
		4504: oled_colour = 16'b00001_000001_00001; 
		4505: oled_colour = 16'b00001_000001_00001; 
		4506: oled_colour = 16'b00001_000001_00001; 
		4507: oled_colour = 16'b00001_000001_00001; 
		4508: oled_colour = 16'b00001_000001_00001; 
		4509: oled_colour = 16'b00001_000001_00001; 
		4510: oled_colour = 16'b00001_000001_00001; 
		4511: oled_colour = 16'b00001_000001_00001; 
		4512: oled_colour = 16'b00001_000001_00001; 
		4513: oled_colour = 16'b00001_000001_00001; 
		4514: oled_colour = 16'b00001_000001_00001; 
		4515: oled_colour = 16'b00001_000001_00001; 
		4516: oled_colour = 16'b00001_000001_00001; 
		4517: oled_colour = 16'b00001_000001_00001; 
		4518: oled_colour = 16'b00001_000001_00001; 
		4519: oled_colour = 16'b00001_000001_00001; 
		4520: oled_colour = 16'b00001_000001_00001; 
		4521: oled_colour = 16'b00001_000001_00001; 
		4522: oled_colour = 16'b00001_000001_00001; 
		4523: oled_colour = 16'b00001_000001_00001; 
		4524: oled_colour = 16'b00001_000001_00001; 
		4525: oled_colour = 16'b00001_000001_00001; 
		4526: oled_colour = 16'b00001_000001_00001; 
		4527: oled_colour = 16'b00001_000001_00001; 
		4528: oled_colour = 16'b00001_000001_00001; 
		4529: oled_colour = 16'b00001_000001_00001; 
		4530: oled_colour = 16'b00001_000001_00001; 
		4531: oled_colour = 16'b00001_000001_00001; 
		4532: oled_colour = 16'b00001_000001_00001; 
		4533: oled_colour = 16'b00001_000001_00001; 
		4534: oled_colour = 16'b00001_000001_00001; 
		4535: oled_colour = 16'b00001_000001_00001; 
		4536: oled_colour = 16'b00001_000001_00001; 
		4537: oled_colour = 16'b00001_000001_00001; 
		4538: oled_colour = 16'b00001_000001_00001; 
		4539: oled_colour = 16'b00001_000001_00001; 
		4540: oled_colour = 16'b00001_000001_00001; 
		4541: oled_colour = 16'b00001_000001_00001; 
		4542: oled_colour = 16'b00001_000001_00001; 
		4543: oled_colour = 16'b00001_000001_00001; 
		4544: oled_colour = 16'b00001_000001_00001; 
		4545: oled_colour = 16'b00001_000001_00001; 
		4546: oled_colour = 16'b00001_000001_00001; 
		4547: oled_colour = 16'b00001_000001_00001; 
		4548: oled_colour = 16'b00001_000001_00001; 
		4549: oled_colour = 16'b00001_000001_00001; 
		4550: oled_colour = 16'b00001_000001_00001; 
		4551: oled_colour = 16'b00001_000001_00001; 
		4552: oled_colour = 16'b00001_000001_00001; 
		4553: oled_colour = 16'b00001_000001_00001; 
		4554: oled_colour = 16'b00001_000001_00001; 
		4555: oled_colour = 16'b00001_000001_00001; 
		4556: oled_colour = 16'b00001_000001_00001; 
		4557: oled_colour = 16'b00001_000001_00001; 
		4558: oled_colour = 16'b00001_000001_00001; 
		4559: oled_colour = 16'b00001_000001_00001; 
		4560: oled_colour = 16'b00001_000001_00001; 
		4561: oled_colour = 16'b00001_000001_00001; 
		4562: oled_colour = 16'b00001_000001_00001; 
		4563: oled_colour = 16'b00001_000001_00001; 
		4564: oled_colour = 16'b00001_000001_00001; 
		4565: oled_colour = 16'b00001_000001_00001; 
		4566: oled_colour = 16'b00001_000001_00001; 
		4567: oled_colour = 16'b00001_000001_00001; 
		4568: oled_colour = 16'b00001_000001_00001; 
		4569: oled_colour = 16'b00001_000001_00001; 
		4570: oled_colour = 16'b00001_000001_00001; 
		4571: oled_colour = 16'b00001_000001_00001; 
		4572: oled_colour = 16'b00001_000001_00001; 
		4573: oled_colour = 16'b00001_000001_00001; 
		4574: oled_colour = 16'b00001_000001_00001; 
		4575: oled_colour = 16'b00001_000001_00001; 
		4576: oled_colour = 16'b00001_000001_00001; 
		4577: oled_colour = 16'b00001_000001_00001; 
		4578: oled_colour = 16'b00001_000001_00001; 
		4579: oled_colour = 16'b00001_000001_00001; 
		4580: oled_colour = 16'b00001_000001_00001; 
		4581: oled_colour = 16'b00001_000001_00001; 
		4582: oled_colour = 16'b00001_000001_00001; 
		4583: oled_colour = 16'b00001_000001_00001; 
		4584: oled_colour = 16'b00001_000001_00001; 
		4585: oled_colour = 16'b00001_000001_00001; 
		4586: oled_colour = 16'b00001_000001_00001; 
		4587: oled_colour = 16'b00001_000001_00001; 
		4588: oled_colour = 16'b00001_000001_00001; 
		4589: oled_colour = 16'b00001_000001_00001; 
		4590: oled_colour = 16'b00001_000001_00001; 
		4591: oled_colour = 16'b00001_000001_00001; 
		4592: oled_colour = 16'b00001_000001_00001; 
		4593: oled_colour = 16'b00001_000001_00001; 
		4594: oled_colour = 16'b00001_000001_00001; 
		4595: oled_colour = 16'b00001_000001_00001; 
		4596: oled_colour = 16'b00001_000001_00001; 
		4597: oled_colour = 16'b00001_000001_00001; 
		4598: oled_colour = 16'b00001_000001_00001; 
		4599: oled_colour = 16'b00001_000001_00001; 
		4600: oled_colour = 16'b00001_000001_00001; 
		4601: oled_colour = 16'b00001_000001_00001; 
		4602: oled_colour = 16'b00001_000001_00001; 
		4603: oled_colour = 16'b00001_000001_00001; 
		4604: oled_colour = 16'b00001_000001_00001; 
		4605: oled_colour = 16'b00001_000001_00001; 
		4606: oled_colour = 16'b00001_000001_00001; 
		4607: oled_colour = 16'b00001_000001_00001; 
		4608: oled_colour = 16'b00001_000001_00001; 
		4609: oled_colour = 16'b00001_000001_00001; 
		4610: oled_colour = 16'b00001_000001_00001; 
		4611: oled_colour = 16'b00001_000001_00001; 
		4612: oled_colour = 16'b00001_000001_00001; 
		4613: oled_colour = 16'b00001_000001_00001; 
		4614: oled_colour = 16'b00001_000001_00001; 
		4615: oled_colour = 16'b00001_000001_00001; 
		4616: oled_colour = 16'b00001_000001_00001; 
		4617: oled_colour = 16'b00001_000001_00001; 
		4618: oled_colour = 16'b00001_000001_00001; 
		4619: oled_colour = 16'b00001_000001_00001; 
		4620: oled_colour = 16'b00001_000001_00001; 
		4621: oled_colour = 16'b00001_000001_00001; 
		4622: oled_colour = 16'b00001_000001_00001; 
		4623: oled_colour = 16'b00001_000001_00001; 
		4624: oled_colour = 16'b00001_000001_00001; 
		4625: oled_colour = 16'b00001_000001_00001; 
		4626: oled_colour = 16'b00001_000001_00001; 
		4627: oled_colour = 16'b00001_000001_00001; 
		4628: oled_colour = 16'b00001_000001_00001; 
		4629: oled_colour = 16'b00001_000001_00001; 
		4630: oled_colour = 16'b00001_000001_00001; 
		4631: oled_colour = 16'b00001_000001_00001; 
		4632: oled_colour = 16'b00001_000001_00001; 
		4633: oled_colour = 16'b00001_000001_00001; 
		4634: oled_colour = 16'b00001_000001_00001; 
		4635: oled_colour = 16'b00001_000001_00001; 
		4636: oled_colour = 16'b00001_000001_00001; 
		4637: oled_colour = 16'b00001_000001_00001; 
		4638: oled_colour = 16'b00001_000001_00001; 
		4639: oled_colour = 16'b00001_000001_00001; 
		4640: oled_colour = 16'b00001_000001_00001; 
		4641: oled_colour = 16'b00001_000001_00001; 
		4642: oled_colour = 16'b00001_000001_00001; 
		4643: oled_colour = 16'b00001_000001_00001; 
		4644: oled_colour = 16'b00001_000001_00001; 
		4645: oled_colour = 16'b00001_000001_00001; 
		4646: oled_colour = 16'b00001_000001_00001; 
		4647: oled_colour = 16'b00001_000001_00001; 
		4648: oled_colour = 16'b00001_000001_00001; 
		4649: oled_colour = 16'b00001_000001_00001; 
		4650: oled_colour = 16'b00001_000001_00001; 
		4651: oled_colour = 16'b00001_000001_00001; 
		4652: oled_colour = 16'b00001_000001_00001; 
		4653: oled_colour = 16'b00001_000001_00001; 
		4654: oled_colour = 16'b00001_000001_00001; 
		4655: oled_colour = 16'b00001_000001_00001; 
		4656: oled_colour = 16'b00001_000001_00001; 
		4657: oled_colour = 16'b00001_000001_00001; 
		4658: oled_colour = 16'b00001_000001_00001; 
		4659: oled_colour = 16'b00001_000001_00001; 
		4660: oled_colour = 16'b00001_000001_00001; 
		4661: oled_colour = 16'b00001_000001_00001; 
		4662: oled_colour = 16'b00001_000001_00001; 
		4663: oled_colour = 16'b00001_000001_00001; 
		4664: oled_colour = 16'b00001_000001_00001; 
		4665: oled_colour = 16'b00001_000001_00001; 
		4666: oled_colour = 16'b00001_000001_00001; 
		4667: oled_colour = 16'b00001_000001_00001; 
		4668: oled_colour = 16'b00001_000001_00001; 
		4669: oled_colour = 16'b00001_000001_00001; 
		4670: oled_colour = 16'b00001_000001_00001; 
		4671: oled_colour = 16'b00001_000001_00001; 
		4672: oled_colour = 16'b00001_000001_00001; 
		4673: oled_colour = 16'b00001_000001_00001; 
		4674: oled_colour = 16'b00001_000001_00001; 
		4675: oled_colour = 16'b00001_000001_00001; 
		4676: oled_colour = 16'b00001_000001_00001; 
		4677: oled_colour = 16'b00001_000001_00001; 
		4678: oled_colour = 16'b00001_000001_00001; 
		4679: oled_colour = 16'b00001_000001_00001; 
		4680: oled_colour = 16'b00001_000001_00001; 
		4681: oled_colour = 16'b00001_000001_00001; 
		4682: oled_colour = 16'b00001_000001_00001; 
		4683: oled_colour = 16'b00001_000001_00001; 
		4684: oled_colour = 16'b00001_000001_00001; 
		4685: oled_colour = 16'b00001_000001_00001; 
		4686: oled_colour = 16'b00001_000001_00001; 
		4687: oled_colour = 16'b00001_000001_00001; 
		4688: oled_colour = 16'b00001_000001_00001; 
		4689: oled_colour = 16'b00001_000001_00001; 
		4690: oled_colour = 16'b00001_000001_00001; 
		4691: oled_colour = 16'b00001_000001_00001; 
		4692: oled_colour = 16'b00001_000001_00001; 
		4693: oled_colour = 16'b00001_000001_00001; 
		4694: oled_colour = 16'b00001_000001_00001; 
		4695: oled_colour = 16'b00001_000001_00001; 
		4696: oled_colour = 16'b00001_000001_00001; 
		4697: oled_colour = 16'b00001_000001_00001; 
		4698: oled_colour = 16'b00001_000001_00001; 
		4699: oled_colour = 16'b00001_000001_00001; 
		4700: oled_colour = 16'b00001_000001_00001; 
		4701: oled_colour = 16'b00001_000001_00001; 
		4702: oled_colour = 16'b00001_000001_00001; 
		4703: oled_colour = 16'b00001_000001_00001; 
		4704: oled_colour = 16'b00001_000001_00001; 
		4705: oled_colour = 16'b00001_000001_00001; 
		4706: oled_colour = 16'b00001_000001_00001; 
		4707: oled_colour = 16'b00001_000001_00001; 
		4708: oled_colour = 16'b00001_000001_00001; 
		4709: oled_colour = 16'b00001_000001_00001; 
		4710: oled_colour = 16'b00001_000001_00001; 
		4711: oled_colour = 16'b00001_000001_00001; 
		4712: oled_colour = 16'b00001_000001_00001; 
		4713: oled_colour = 16'b00001_000001_00001; 
		4714: oled_colour = 16'b00001_000001_00001; 
		4715: oled_colour = 16'b00001_000001_00001; 
		4716: oled_colour = 16'b00001_000001_00001; 
		4717: oled_colour = 16'b00001_000001_00001; 
		4718: oled_colour = 16'b00001_000001_00001; 
		4719: oled_colour = 16'b00001_000001_00001; 
		4720: oled_colour = 16'b00001_000001_00001; 
		4721: oled_colour = 16'b00001_000001_00001; 
		4722: oled_colour = 16'b00001_000001_00001; 
		4723: oled_colour = 16'b00001_000001_00001; 
		4724: oled_colour = 16'b00001_000001_00001; 
		4725: oled_colour = 16'b00001_000001_00001; 
		4726: oled_colour = 16'b00001_000001_00001; 
		4727: oled_colour = 16'b00001_000001_00001; 
		4728: oled_colour = 16'b00001_000001_00001; 
		4729: oled_colour = 16'b00001_000001_00001; 
		4730: oled_colour = 16'b00001_000001_00001; 
		4731: oled_colour = 16'b00001_000001_00001; 
		4732: oled_colour = 16'b00001_000001_00001; 
		4733: oled_colour = 16'b00001_000001_00001; 
		4734: oled_colour = 16'b00001_000001_00001; 
		4735: oled_colour = 16'b00001_000001_00001; 
		4736: oled_colour = 16'b00001_000001_00001; 
		4737: oled_colour = 16'b00001_000001_00001; 
		4738: oled_colour = 16'b00001_000001_00001; 
		4739: oled_colour = 16'b00001_000001_00001; 
		4740: oled_colour = 16'b00001_000001_00001; 
		4741: oled_colour = 16'b00001_000001_00001; 
		4742: oled_colour = 16'b00001_000001_00001; 
		4743: oled_colour = 16'b00001_000001_00001; 
		4744: oled_colour = 16'b00001_000001_00001; 
		4745: oled_colour = 16'b00001_000001_00001; 
		4746: oled_colour = 16'b00001_000001_00001; 
		4747: oled_colour = 16'b00001_000001_00001; 
		4748: oled_colour = 16'b00001_000001_00001; 
		4749: oled_colour = 16'b00001_000001_00001; 
		4750: oled_colour = 16'b00001_000001_00001; 
		4751: oled_colour = 16'b00001_000001_00001; 
		4752: oled_colour = 16'b00001_000001_00001; 
		4753: oled_colour = 16'b00001_000001_00001; 
		4754: oled_colour = 16'b00001_000001_00001; 
		4755: oled_colour = 16'b00001_000001_00001; 
		4756: oled_colour = 16'b00001_000001_00001; 
		4757: oled_colour = 16'b00001_000001_00001; 
		4758: oled_colour = 16'b00001_000001_00001; 
		4759: oled_colour = 16'b00001_000001_00001; 
		4760: oled_colour = 16'b00001_000001_00001; 
		4761: oled_colour = 16'b00001_000001_00001; 
		4762: oled_colour = 16'b00001_000001_00001; 
		4763: oled_colour = 16'b00001_000001_00001; 
		4764: oled_colour = 16'b00001_000001_00001; 
		4765: oled_colour = 16'b00001_000001_00001; 
		4766: oled_colour = 16'b00001_000001_00001; 
		4767: oled_colour = 16'b00001_000001_00001; 
		4768: oled_colour = 16'b00001_000001_00001; 
		4769: oled_colour = 16'b00001_000001_00001; 
		4770: oled_colour = 16'b00001_000001_00001; 
		4771: oled_colour = 16'b00001_000001_00001; 
		4772: oled_colour = 16'b00001_000001_00001; 
		4773: oled_colour = 16'b00001_000001_00001; 
		4774: oled_colour = 16'b00001_000001_00001; 
		4775: oled_colour = 16'b00001_000001_00001; 
		4776: oled_colour = 16'b00001_000001_00001; 
		4777: oled_colour = 16'b00001_000001_00001; 
		4778: oled_colour = 16'b00001_000001_00001; 
		4779: oled_colour = 16'b00001_000001_00001; 
		4780: oled_colour = 16'b00001_000001_00001; 
		4781: oled_colour = 16'b00001_000001_00001; 
		4782: oled_colour = 16'b00001_000001_00001; 
		4783: oled_colour = 16'b00001_000001_00001; 
		4784: oled_colour = 16'b00001_000001_00001; 
		4785: oled_colour = 16'b00001_000001_00001; 
		4786: oled_colour = 16'b00001_000001_00001; 
		4787: oled_colour = 16'b00001_000001_00001; 
		4788: oled_colour = 16'b00001_000001_00001; 
		4789: oled_colour = 16'b00001_000001_00001; 
		4790: oled_colour = 16'b00001_000001_00001; 
		4791: oled_colour = 16'b00001_000001_00001; 
		4792: oled_colour = 16'b00001_000001_00001; 
		4793: oled_colour = 16'b00001_000001_00001; 
		4794: oled_colour = 16'b00001_000001_00001; 
		4795: oled_colour = 16'b00001_000001_00001; 
		4796: oled_colour = 16'b00001_000001_00001; 
		4797: oled_colour = 16'b00001_000001_00001; 
		4798: oled_colour = 16'b00001_000001_00001; 
		4799: oled_colour = 16'b00001_000001_00001; 
		4800: oled_colour = 16'b00001_000001_00001; 
		4801: oled_colour = 16'b00001_000001_00001; 
		4802: oled_colour = 16'b00001_000001_00001; 
		4803: oled_colour = 16'b00001_000001_00001; 
		4804: oled_colour = 16'b00001_000001_00001; 
		4805: oled_colour = 16'b00001_000001_00001; 
		4806: oled_colour = 16'b00001_000001_00001; 
		4807: oled_colour = 16'b00001_000001_00001; 
		4808: oled_colour = 16'b00001_000001_00001; 
		4809: oled_colour = 16'b00001_000001_00001; 
		4810: oled_colour = 16'b00001_000001_00001; 
		4811: oled_colour = 16'b00001_000001_00001; 
		4812: oled_colour = 16'b00001_000001_00001; 
		4813: oled_colour = 16'b00001_000001_00001; 
		4814: oled_colour = 16'b00001_000001_00001; 
		4815: oled_colour = 16'b00001_000001_00001; 
		4816: oled_colour = 16'b00001_000001_00001; 
		4817: oled_colour = 16'b00001_000001_00001; 
		4818: oled_colour = 16'b00001_000001_00001; 
		4819: oled_colour = 16'b00001_000001_00001; 
		4820: oled_colour = 16'b00001_000001_00001; 
		4821: oled_colour = 16'b00001_000001_00001; 
		4822: oled_colour = 16'b00001_000001_00001; 
		4823: oled_colour = 16'b00001_000001_00001; 
		4824: oled_colour = 16'b00001_000001_00001; 
		4825: oled_colour = 16'b00001_000001_00001; 
		4826: oled_colour = 16'b00001_000001_00001; 
		4827: oled_colour = 16'b00001_000001_00001; 
		4828: oled_colour = 16'b00001_000001_00001; 
		4829: oled_colour = 16'b00001_000001_00001; 
		4830: oled_colour = 16'b00001_000001_00001; 
		4831: oled_colour = 16'b00001_000001_00001; 
		4832: oled_colour = 16'b00001_000001_00001; 
		4833: oled_colour = 16'b00001_000001_00001; 
		4834: oled_colour = 16'b00001_000001_00001; 
		4835: oled_colour = 16'b00001_000001_00001; 
		4836: oled_colour = 16'b00001_000001_00001; 
		4837: oled_colour = 16'b00001_000001_00001; 
		4838: oled_colour = 16'b00001_000001_00001; 
		4839: oled_colour = 16'b00001_000001_00001; 
		4840: oled_colour = 16'b00001_000001_00001; 
		4841: oled_colour = 16'b00001_000001_00001; 
		4842: oled_colour = 16'b00001_000001_00001; 
		4843: oled_colour = 16'b00001_000001_00001; 
		4844: oled_colour = 16'b00001_000001_00001; 
		4845: oled_colour = 16'b00001_000001_00001; 
		4846: oled_colour = 16'b00001_000001_00001; 
		4847: oled_colour = 16'b00001_000001_00001; 
		4848: oled_colour = 16'b00001_000001_00001; 
		4849: oled_colour = 16'b00001_000001_00001; 
		4850: oled_colour = 16'b00001_000001_00001; 
		4851: oled_colour = 16'b00001_000001_00001; 
		4852: oled_colour = 16'b00001_000001_00001; 
		4853: oled_colour = 16'b00001_000001_00001; 
		4854: oled_colour = 16'b00001_000001_00001; 
		4855: oled_colour = 16'b00001_000001_00001; 
		4856: oled_colour = 16'b00001_000001_00001; 
		4857: oled_colour = 16'b00001_000001_00001; 
		4858: oled_colour = 16'b00001_000001_00001; 
		4859: oled_colour = 16'b00001_000001_00001; 
		4860: oled_colour = 16'b00001_000001_00001; 
		4861: oled_colour = 16'b00001_000001_00001; 
		4862: oled_colour = 16'b00001_000001_00001; 
		4863: oled_colour = 16'b00001_000001_00001; 
		4864: oled_colour = 16'b00001_000001_00001; 
		4865: oled_colour = 16'b00001_000001_00001; 
		4866: oled_colour = 16'b00001_000001_00001; 
		4867: oled_colour = 16'b00001_000001_00001; 
		4868: oled_colour = 16'b00001_000001_00001; 
		4869: oled_colour = 16'b00001_000001_00001; 
		4870: oled_colour = 16'b00001_000001_00001; 
		4871: oled_colour = 16'b00001_000001_00001; 
		4872: oled_colour = 16'b00001_000001_00001; 
		4873: oled_colour = 16'b00001_000001_00001; 
		4874: oled_colour = 16'b00001_000001_00001; 
		4875: oled_colour = 16'b00001_000001_00001; 
		4876: oled_colour = 16'b00001_000001_00001; 
		4877: oled_colour = 16'b00001_000001_00001; 
		4878: oled_colour = 16'b00001_000001_00001; 
		4879: oled_colour = 16'b00001_000001_00001; 
		4880: oled_colour = 16'b00001_000001_00001; 
		4881: oled_colour = 16'b00001_000001_00001; 
		4882: oled_colour = 16'b00001_000001_00001; 
		4883: oled_colour = 16'b00001_000001_00001; 
		4884: oled_colour = 16'b00001_000001_00001; 
		4885: oled_colour = 16'b00001_000001_00001; 
		4886: oled_colour = 16'b00001_000001_00001; 
		4887: oled_colour = 16'b00001_000001_00001; 
		4888: oled_colour = 16'b00001_000001_00001; 
		4889: oled_colour = 16'b00001_000001_00001; 
		4890: oled_colour = 16'b00001_000001_00001; 
		4891: oled_colour = 16'b00001_000001_00001; 
		4892: oled_colour = 16'b00001_000001_00001; 
		4893: oled_colour = 16'b00001_000001_00001; 
		4894: oled_colour = 16'b00001_000001_00001; 
		4895: oled_colour = 16'b00001_000001_00001; 
		4896: oled_colour = 16'b00001_000001_00001; 
		4897: oled_colour = 16'b00001_000001_00001; 
		4898: oled_colour = 16'b00001_000001_00001; 
		4899: oled_colour = 16'b00001_000001_00001; 
		4900: oled_colour = 16'b00001_000001_00001; 
		4901: oled_colour = 16'b00001_000001_00001; 
		4902: oled_colour = 16'b00001_000001_00001; 
		4903: oled_colour = 16'b00001_000001_00001; 
		4904: oled_colour = 16'b00001_000001_00001; 
		4905: oled_colour = 16'b00001_000001_00001; 
		4906: oled_colour = 16'b00001_000001_00001; 
		4907: oled_colour = 16'b00001_000001_00001; 
		4908: oled_colour = 16'b00001_000001_00001; 
		4909: oled_colour = 16'b00001_000001_00001; 
		4910: oled_colour = 16'b00001_000001_00001; 
		4911: oled_colour = 16'b00001_000001_00001; 
		4912: oled_colour = 16'b00001_000001_00001; 
		4913: oled_colour = 16'b00001_000001_00001; 
		4914: oled_colour = 16'b00001_000001_00001; 
		4915: oled_colour = 16'b00001_000001_00001; 
		4916: oled_colour = 16'b00001_000001_00001; 
		4917: oled_colour = 16'b00001_000001_00001; 
		4918: oled_colour = 16'b00001_000001_00001; 
		4919: oled_colour = 16'b00001_000001_00001; 
		4920: oled_colour = 16'b00001_000001_00001; 
		4921: oled_colour = 16'b00001_000001_00001; 
		4922: oled_colour = 16'b00001_000001_00001; 
		4923: oled_colour = 16'b00001_000001_00001; 
		4924: oled_colour = 16'b00001_000001_00001; 
		4925: oled_colour = 16'b00001_000001_00001; 
		4926: oled_colour = 16'b00001_000001_00001; 
		4927: oled_colour = 16'b00001_000001_00001; 
		4928: oled_colour = 16'b00001_000001_00001; 
		4929: oled_colour = 16'b00001_000001_00001; 
		4930: oled_colour = 16'b00001_000001_00001; 
		4931: oled_colour = 16'b00001_000001_00001; 
		4932: oled_colour = 16'b00001_000001_00001; 
		4933: oled_colour = 16'b00001_000001_00001; 
		4934: oled_colour = 16'b00001_000001_00001; 
		4935: oled_colour = 16'b00001_000001_00001; 
		4936: oled_colour = 16'b00001_000001_00001; 
		4937: oled_colour = 16'b00001_000001_00001; 
		4938: oled_colour = 16'b00001_000001_00001; 
		4939: oled_colour = 16'b00001_000001_00001; 
		4940: oled_colour = 16'b00001_000001_00001; 
		4941: oled_colour = 16'b00001_000001_00001; 
		4942: oled_colour = 16'b00001_000001_00001; 
		4943: oled_colour = 16'b00001_000001_00001; 
		4944: oled_colour = 16'b00001_000001_00001; 
		4945: oled_colour = 16'b00001_000001_00001; 
		4946: oled_colour = 16'b00001_000001_00001; 
		4947: oled_colour = 16'b00001_000001_00001; 
		4948: oled_colour = 16'b00001_000001_00001; 
		4949: oled_colour = 16'b00001_000001_00001; 
		4950: oled_colour = 16'b00001_000001_00001; 
		4951: oled_colour = 16'b00001_000001_00001; 
		4952: oled_colour = 16'b00001_000001_00001; 
		4953: oled_colour = 16'b00001_000001_00001; 
		4954: oled_colour = 16'b00001_000001_00001; 
		4955: oled_colour = 16'b00001_000001_00001; 
		4956: oled_colour = 16'b00001_000001_00001; 
		4957: oled_colour = 16'b00001_000001_00001; 
		4958: oled_colour = 16'b00001_000001_00001; 
		4959: oled_colour = 16'b00001_000001_00001; 
		4960: oled_colour = 16'b00001_000001_00001; 
		4961: oled_colour = 16'b00001_000001_00001; 
		4962: oled_colour = 16'b00001_000001_00001; 
		4963: oled_colour = 16'b00001_000001_00001; 
		4964: oled_colour = 16'b00001_000001_00001; 
		4965: oled_colour = 16'b00001_000001_00001; 
		4966: oled_colour = 16'b00001_000001_00001; 
		4967: oled_colour = 16'b00001_000001_00001; 
		4968: oled_colour = 16'b00001_000001_00001; 
		4969: oled_colour = 16'b00001_000001_00001; 
		4970: oled_colour = 16'b00001_000001_00001; 
		4971: oled_colour = 16'b00001_000001_00001; 
		4972: oled_colour = 16'b00001_000001_00001; 
		4973: oled_colour = 16'b00001_000001_00001; 
		4974: oled_colour = 16'b00001_000001_00001; 
		4975: oled_colour = 16'b00001_000001_00001; 
		4976: oled_colour = 16'b00001_000001_00001; 
		4977: oled_colour = 16'b00001_000001_00001; 
		4978: oled_colour = 16'b00001_000001_00001; 
		4979: oled_colour = 16'b00001_000001_00001; 
		4980: oled_colour = 16'b00001_000001_00001; 
		4981: oled_colour = 16'b00001_000001_00001; 
		4982: oled_colour = 16'b00001_000001_00001; 
		4983: oled_colour = 16'b00001_000001_00001; 
		4984: oled_colour = 16'b00001_000001_00001; 
		4985: oled_colour = 16'b00001_000001_00001; 
		4986: oled_colour = 16'b00001_000001_00001; 
		4987: oled_colour = 16'b00001_000001_00001; 
		4988: oled_colour = 16'b00001_000001_00001; 
		4989: oled_colour = 16'b00001_000001_00001; 
		4990: oled_colour = 16'b00001_000001_00001; 
		4991: oled_colour = 16'b00001_000001_00001; 
		4992: oled_colour = 16'b00001_000001_00001; 
		4993: oled_colour = 16'b00001_000001_00001; 
		4994: oled_colour = 16'b00001_000001_00001; 
		4995: oled_colour = 16'b00001_000001_00001; 
		4996: oled_colour = 16'b00001_000001_00001; 
		4997: oled_colour = 16'b00001_000001_00001; 
		4998: oled_colour = 16'b00001_000001_00001; 
		4999: oled_colour = 16'b00001_000001_00001; 
		5000: oled_colour = 16'b00001_000001_00001; 
		5001: oled_colour = 16'b00001_000001_00001; 
		5002: oled_colour = 16'b00001_000001_00001; 
		5003: oled_colour = 16'b00001_000001_00001; 
		5004: oled_colour = 16'b00001_000001_00001; 
		5005: oled_colour = 16'b00001_000001_00001; 
		5006: oled_colour = 16'b00001_000001_00001; 
		5007: oled_colour = 16'b00001_000001_00001; 
		5008: oled_colour = 16'b00001_000001_00001; 
		5009: oled_colour = 16'b00001_000001_00001; 
		5010: oled_colour = 16'b00001_000001_00001; 
		5011: oled_colour = 16'b00001_000001_00001; 
		5012: oled_colour = 16'b00001_000001_00001; 
		5013: oled_colour = 16'b00001_000001_00001; 
		5014: oled_colour = 16'b00001_000001_00001; 
		5015: oled_colour = 16'b00001_000001_00001; 
		5016: oled_colour = 16'b00001_000001_00001; 
		5017: oled_colour = 16'b00001_000001_00001; 
		5018: oled_colour = 16'b00001_000001_00001; 
		5019: oled_colour = 16'b00001_000001_00001; 
		5020: oled_colour = 16'b00001_000001_00001; 
		5021: oled_colour = 16'b00001_000001_00001; 
		5022: oled_colour = 16'b00001_000001_00001; 
		5023: oled_colour = 16'b00001_000001_00001; 
		5024: oled_colour = 16'b00001_000001_00001; 
		5025: oled_colour = 16'b00001_000001_00001; 
		5026: oled_colour = 16'b00001_000001_00001; 
		5027: oled_colour = 16'b00001_000001_00001; 
		5028: oled_colour = 16'b00001_000001_00001; 
		5029: oled_colour = 16'b00001_000001_00001; 
		5030: oled_colour = 16'b00001_000001_00001; 
		5031: oled_colour = 16'b00001_000001_00001; 
		5032: oled_colour = 16'b00001_000001_00001; 
		5033: oled_colour = 16'b00001_000001_00001; 
		5034: oled_colour = 16'b00001_000001_00001; 
		5035: oled_colour = 16'b00001_000001_00001; 
		5036: oled_colour = 16'b00001_000001_00001; 
		5037: oled_colour = 16'b00001_000001_00001; 
		5038: oled_colour = 16'b00001_000001_00001; 
		5039: oled_colour = 16'b00001_000001_00001; 
		5040: oled_colour = 16'b00001_000001_00001; 
		5041: oled_colour = 16'b00001_000001_00001; 
		5042: oled_colour = 16'b00001_000001_00001; 
		5043: oled_colour = 16'b00001_000001_00001; 
		5044: oled_colour = 16'b00001_000001_00001; 
		5045: oled_colour = 16'b00001_000001_00001; 
		5046: oled_colour = 16'b00001_000001_00001; 
		5047: oled_colour = 16'b00001_000001_00001; 
		5048: oled_colour = 16'b00001_000001_00001; 
		5049: oled_colour = 16'b00001_000001_00001; 
		5050: oled_colour = 16'b00001_000001_00001; 
		5051: oled_colour = 16'b00001_000001_00001; 
		5052: oled_colour = 16'b00001_000001_00001; 
		5053: oled_colour = 16'b00001_000001_00001; 
		5054: oled_colour = 16'b00001_000001_00001; 
		5055: oled_colour = 16'b00001_000001_00001; 
		5056: oled_colour = 16'b00001_000001_00001; 
		5057: oled_colour = 16'b00001_000001_00001; 
		5058: oled_colour = 16'b00001_000001_00001; 
		5059: oled_colour = 16'b00001_000001_00001; 
		5060: oled_colour = 16'b00001_000001_00001; 
		5061: oled_colour = 16'b00001_000001_00001; 
		5062: oled_colour = 16'b00001_000001_00001; 
		5063: oled_colour = 16'b00001_000001_00001; 
		5064: oled_colour = 16'b00001_000001_00001; 
		5065: oled_colour = 16'b00001_000001_00001; 
		5066: oled_colour = 16'b00001_000001_00001; 
		5067: oled_colour = 16'b00001_000001_00001; 
		5068: oled_colour = 16'b00001_000001_00001; 
		5069: oled_colour = 16'b00001_000001_00001; 
		5070: oled_colour = 16'b00001_000001_00001; 
		5071: oled_colour = 16'b00001_000001_00001; 
		5072: oled_colour = 16'b00001_000001_00001; 
		5073: oled_colour = 16'b00001_000001_00001; 
		5074: oled_colour = 16'b00001_000001_00001; 
		5075: oled_colour = 16'b00001_000001_00001; 
		5076: oled_colour = 16'b00001_000001_00001; 
		5077: oled_colour = 16'b00001_000001_00001; 
		5078: oled_colour = 16'b00001_000001_00001; 
		5079: oled_colour = 16'b00001_000001_00001; 
		5080: oled_colour = 16'b00001_000001_00001; 
		5081: oled_colour = 16'b00001_000001_00001; 
		5082: oled_colour = 16'b00001_000001_00001; 
		5083: oled_colour = 16'b00001_000001_00001; 
		5084: oled_colour = 16'b00001_000001_00001; 
		5085: oled_colour = 16'b00001_000001_00001; 
		5086: oled_colour = 16'b00001_000001_00001; 
		5087: oled_colour = 16'b00001_000001_00001; 
		5088: oled_colour = 16'b00001_000001_00001; 
		5089: oled_colour = 16'b00001_000001_00001; 
		5090: oled_colour = 16'b00001_000001_00001; 
		5091: oled_colour = 16'b00001_000001_00001; 
		5092: oled_colour = 16'b00001_000001_00001; 
		5093: oled_colour = 16'b00001_000001_00001; 
		5094: oled_colour = 16'b00001_000001_00001; 
		5095: oled_colour = 16'b00001_000001_00001; 
		5096: oled_colour = 16'b00001_000001_00001; 
		5097: oled_colour = 16'b00001_000001_00001; 
		5098: oled_colour = 16'b00001_000001_00001; 
		5099: oled_colour = 16'b00001_000001_00001; 
		5100: oled_colour = 16'b00001_000001_00001; 
		5101: oled_colour = 16'b00001_000001_00001; 
		5102: oled_colour = 16'b00001_000001_00001; 
		5103: oled_colour = 16'b00001_000001_00001; 
		5104: oled_colour = 16'b00001_000001_00001; 
		5105: oled_colour = 16'b00001_000001_00001; 
		5106: oled_colour = 16'b00001_000001_00001; 
		5107: oled_colour = 16'b00001_000001_00001; 
		5108: oled_colour = 16'b00001_000001_00001; 
		5109: oled_colour = 16'b00001_000001_00001; 
		5110: oled_colour = 16'b00001_000001_00001; 
		5111: oled_colour = 16'b00001_000001_00001; 
		5112: oled_colour = 16'b00001_000001_00001; 
		5113: oled_colour = 16'b00001_000001_00001; 
		5114: oled_colour = 16'b00001_000001_00001; 
		5115: oled_colour = 16'b00001_000001_00001; 
		5116: oled_colour = 16'b00001_000001_00001; 
		5117: oled_colour = 16'b00001_000001_00001; 
		5118: oled_colour = 16'b00001_000001_00001; 
		5119: oled_colour = 16'b00001_000001_00001; 
		5120: oled_colour = 16'b00001_000001_00001; 
		5121: oled_colour = 16'b00001_000001_00001; 
		5122: oled_colour = 16'b00001_000001_00001; 
		5123: oled_colour = 16'b00001_000001_00001; 
		5124: oled_colour = 16'b00001_000001_00001; 
		5125: oled_colour = 16'b00001_000001_00001; 
		5126: oled_colour = 16'b00001_000001_00001; 
		5127: oled_colour = 16'b00001_000001_00001; 
		5128: oled_colour = 16'b00001_000001_00001; 
		5129: oled_colour = 16'b00001_000001_00001; 
		5130: oled_colour = 16'b00001_000001_00001; 
		5131: oled_colour = 16'b00001_000001_00001; 
		5132: oled_colour = 16'b00001_000001_00001; 
		5133: oled_colour = 16'b00001_000001_00001; 
		5134: oled_colour = 16'b00001_000001_00001; 
		5135: oled_colour = 16'b00001_000001_00001; 
		5136: oled_colour = 16'b00001_000001_00001; 
		5137: oled_colour = 16'b00001_000001_00001; 
		5138: oled_colour = 16'b00001_000001_00001; 
		5139: oled_colour = 16'b00001_000001_00001; 
		5140: oled_colour = 16'b00001_000001_00001; 
		5141: oled_colour = 16'b00001_000001_00001; 
		5142: oled_colour = 16'b00001_000001_00001; 
		5143: oled_colour = 16'b00001_000001_00001; 
		5144: oled_colour = 16'b00001_000001_00001; 
		5145: oled_colour = 16'b00001_000001_00001; 
		5146: oled_colour = 16'b00001_000001_00001; 
		5147: oled_colour = 16'b00001_000001_00001; 
		5148: oled_colour = 16'b00001_000001_00001; 
		5149: oled_colour = 16'b00001_000001_00001; 
		5150: oled_colour = 16'b00001_000001_00001; 
		5151: oled_colour = 16'b00001_000001_00001; 
		5152: oled_colour = 16'b00001_000001_00001; 
		5153: oled_colour = 16'b00001_000001_00001; 
		5154: oled_colour = 16'b00001_000001_00001; 
		5155: oled_colour = 16'b00001_000001_00001; 
		5156: oled_colour = 16'b00001_000001_00001; 
		5157: oled_colour = 16'b00001_000001_00001; 
		5158: oled_colour = 16'b00001_000001_00001; 
		5159: oled_colour = 16'b00001_000001_00001; 
		5160: oled_colour = 16'b00001_000001_00001; 
		5161: oled_colour = 16'b00001_000001_00001; 
		5162: oled_colour = 16'b00001_000001_00001; 
		5163: oled_colour = 16'b00001_000001_00001; 
		5164: oled_colour = 16'b00001_000001_00001; 
		5165: oled_colour = 16'b00001_000001_00001; 
		5166: oled_colour = 16'b00001_000001_00001; 
		5167: oled_colour = 16'b00001_000001_00001; 
		5168: oled_colour = 16'b00001_000001_00001; 
		5169: oled_colour = 16'b00001_000001_00001; 
		5170: oled_colour = 16'b00001_000001_00001; 
		5171: oled_colour = 16'b00001_000001_00001; 
		5172: oled_colour = 16'b00001_000001_00001; 
		5173: oled_colour = 16'b00001_000001_00001; 
		5174: oled_colour = 16'b00001_000001_00001; 
		5175: oled_colour = 16'b00001_000001_00001; 
		5176: oled_colour = 16'b00001_000001_00001; 
		5177: oled_colour = 16'b00001_000001_00001; 
		5178: oled_colour = 16'b00001_000001_00001; 
		5179: oled_colour = 16'b00001_000001_00001; 
		5180: oled_colour = 16'b00001_000001_00001; 
		5181: oled_colour = 16'b00001_000001_00001; 
		5182: oled_colour = 16'b00001_000001_00001; 
		5183: oled_colour = 16'b00001_000001_00001; 
		5184: oled_colour = 16'b00001_000001_00001; 
		5185: oled_colour = 16'b00001_000001_00001; 
		5186: oled_colour = 16'b00001_000001_00001; 
		5187: oled_colour = 16'b00001_000001_00001; 
		5188: oled_colour = 16'b00001_000001_00001; 
		5189: oled_colour = 16'b00001_000001_00001; 
		5190: oled_colour = 16'b00001_000001_00001; 
		5191: oled_colour = 16'b00001_000001_00001; 
		5192: oled_colour = 16'b00001_000001_00001; 
		5193: oled_colour = 16'b00001_000001_00001; 
		5194: oled_colour = 16'b00001_000001_00001; 
		5195: oled_colour = 16'b00001_000001_00001; 
		5196: oled_colour = 16'b00001_000001_00001; 
		5197: oled_colour = 16'b00001_000001_00001; 
		5198: oled_colour = 16'b00001_000001_00001; 
		5199: oled_colour = 16'b00001_000001_00001; 
		5200: oled_colour = 16'b00001_000001_00001; 
		5201: oled_colour = 16'b00001_000001_00001; 
		5202: oled_colour = 16'b00001_000001_00001; 
		5203: oled_colour = 16'b00001_000001_00001; 
		5204: oled_colour = 16'b00001_000001_00001; 
		5205: oled_colour = 16'b00001_000001_00001; 
		5206: oled_colour = 16'b00001_000001_00001; 
		5207: oled_colour = 16'b00001_000001_00001; 
		5208: oled_colour = 16'b00001_000001_00001; 
		5209: oled_colour = 16'b00001_000001_00001; 
		5210: oled_colour = 16'b00001_000001_00001; 
		5211: oled_colour = 16'b00001_000001_00001; 
		5212: oled_colour = 16'b00001_000001_00001; 
		5213: oled_colour = 16'b00001_000001_00001; 
		5214: oled_colour = 16'b00001_000001_00001; 
		5215: oled_colour = 16'b00001_000001_00001; 
		5216: oled_colour = 16'b00001_000001_00001; 
		5217: oled_colour = 16'b00001_000001_00001; 
		5218: oled_colour = 16'b00001_000001_00001; 
		5219: oled_colour = 16'b00001_000001_00001; 
		5220: oled_colour = 16'b00001_000001_00001; 
		5221: oled_colour = 16'b00001_000001_00001; 
		5222: oled_colour = 16'b00001_000001_00001; 
		5223: oled_colour = 16'b00001_000001_00001; 
		5224: oled_colour = 16'b00001_000001_00001; 
		5225: oled_colour = 16'b00001_000001_00001; 
		5226: oled_colour = 16'b00001_000001_00001; 
		5227: oled_colour = 16'b00001_000001_00001; 
		5228: oled_colour = 16'b00001_000001_00001; 
		5229: oled_colour = 16'b00001_000001_00001; 
		5230: oled_colour = 16'b00001_000001_00001; 
		5231: oled_colour = 16'b00001_000001_00001; 
		5232: oled_colour = 16'b00001_000001_00001; 
		5233: oled_colour = 16'b00001_000001_00001; 
		5234: oled_colour = 16'b00001_000001_00001; 
		5235: oled_colour = 16'b00001_000001_00001; 
		5236: oled_colour = 16'b00001_000001_00001; 
		5237: oled_colour = 16'b00001_000001_00001; 
		5238: oled_colour = 16'b00001_000001_00001; 
		5239: oled_colour = 16'b00001_000001_00001; 
		5240: oled_colour = 16'b00001_000001_00001; 
		5241: oled_colour = 16'b00001_000001_00001; 
		5242: oled_colour = 16'b00001_000001_00001; 
		5243: oled_colour = 16'b00001_000001_00001; 
		5244: oled_colour = 16'b00001_000001_00001; 
		5245: oled_colour = 16'b00001_000001_00001; 
		5246: oled_colour = 16'b00001_000001_00001; 
		5247: oled_colour = 16'b00001_000001_00001; 
		5248: oled_colour = 16'b00001_000001_00001; 
		5249: oled_colour = 16'b00001_000001_00001; 
		5250: oled_colour = 16'b00001_000001_00001; 
		5251: oled_colour = 16'b00001_000001_00001; 
		5252: oled_colour = 16'b00001_000001_00001; 
		5253: oled_colour = 16'b00001_000001_00001; 
		5254: oled_colour = 16'b00001_000001_00001; 
		5255: oled_colour = 16'b00001_000001_00001; 
		5256: oled_colour = 16'b00001_000001_00001; 
		5257: oled_colour = 16'b00001_000001_00001; 
		5258: oled_colour = 16'b00001_000001_00001; 
		5259: oled_colour = 16'b00001_000001_00001; 
		5260: oled_colour = 16'b00001_000001_00001; 
		5261: oled_colour = 16'b00001_000001_00001; 
		5262: oled_colour = 16'b00001_000001_00001; 
		5263: oled_colour = 16'b00001_000001_00001; 
		5264: oled_colour = 16'b00001_000001_00001; 
		5265: oled_colour = 16'b00001_000001_00001; 
		5266: oled_colour = 16'b00001_000001_00001; 
		5267: oled_colour = 16'b00001_000001_00001; 
		5268: oled_colour = 16'b00001_000001_00001; 
		5269: oled_colour = 16'b00001_000001_00001; 
		5270: oled_colour = 16'b00001_000001_00001; 
		5271: oled_colour = 16'b00001_000001_00001; 
		5272: oled_colour = 16'b00001_000001_00001; 
		5273: oled_colour = 16'b00001_000001_00001; 
		5274: oled_colour = 16'b00001_000001_00001; 
		5275: oled_colour = 16'b00001_000001_00001; 
		5276: oled_colour = 16'b00001_000001_00001; 
		5277: oled_colour = 16'b00001_000001_00001; 
		5278: oled_colour = 16'b00001_000001_00001; 
		5279: oled_colour = 16'b00001_000001_00001; 
		5280: oled_colour = 16'b00001_000001_00001; 
		5281: oled_colour = 16'b00001_000001_00001; 
		5282: oled_colour = 16'b00001_000001_00001; 
		5283: oled_colour = 16'b00001_000001_00001; 
		5284: oled_colour = 16'b00001_000001_00001; 
		5285: oled_colour = 16'b00001_000001_00001; 
		5286: oled_colour = 16'b00001_000001_00001; 
		5287: oled_colour = 16'b00001_000001_00001; 
		5288: oled_colour = 16'b00001_000001_00001; 
		5289: oled_colour = 16'b00001_000001_00001; 
		5290: oled_colour = 16'b00001_000001_00001; 
		5291: oled_colour = 16'b00001_000001_00001; 
		5292: oled_colour = 16'b00001_000001_00001; 
		5293: oled_colour = 16'b00001_000001_00001; 
		5294: oled_colour = 16'b00001_000001_00001; 
		5295: oled_colour = 16'b00001_000001_00001; 
		5296: oled_colour = 16'b00001_000001_00001; 
		5297: oled_colour = 16'b00001_000001_00001; 
		5298: oled_colour = 16'b00001_000001_00001; 
		5299: oled_colour = 16'b00001_000001_00001; 
		5300: oled_colour = 16'b00001_000001_00001; 
		5301: oled_colour = 16'b00001_000001_00001; 
		5302: oled_colour = 16'b00001_000001_00001; 
		5303: oled_colour = 16'b00001_000001_00001; 
		5304: oled_colour = 16'b00001_000001_00001; 
		5305: oled_colour = 16'b00001_000001_00001; 
		5306: oled_colour = 16'b00001_000001_00001; 
		5307: oled_colour = 16'b00001_000001_00001; 
		5308: oled_colour = 16'b00001_000001_00001; 
		5309: oled_colour = 16'b00001_000001_00001; 
		5310: oled_colour = 16'b00001_000001_00001; 
		5311: oled_colour = 16'b00001_000001_00001; 
		5312: oled_colour = 16'b00001_000001_00001; 
		5313: oled_colour = 16'b00001_000001_00001; 
		5314: oled_colour = 16'b00001_000001_00001; 
		5315: oled_colour = 16'b00001_000001_00001; 
		5316: oled_colour = 16'b00001_000001_00001; 
		5317: oled_colour = 16'b00001_000001_00001; 
		5318: oled_colour = 16'b00001_000001_00001; 
		5319: oled_colour = 16'b00001_000001_00001; 
		5320: oled_colour = 16'b00001_000001_00001; 
		5321: oled_colour = 16'b00001_000001_00001; 
		5322: oled_colour = 16'b00001_000001_00001; 
		5323: oled_colour = 16'b00001_000001_00001; 
		5324: oled_colour = 16'b00001_000001_00001; 
		5325: oled_colour = 16'b00001_000001_00001; 
		5326: oled_colour = 16'b00001_000001_00001; 
		5327: oled_colour = 16'b00001_000001_00001; 
		5328: oled_colour = 16'b00001_000001_00001; 
		5329: oled_colour = 16'b00001_000001_00001; 
		5330: oled_colour = 16'b00001_000001_00001; 
		5331: oled_colour = 16'b00001_000001_00001; 
		5332: oled_colour = 16'b00001_000001_00001; 
		5333: oled_colour = 16'b00001_000001_00001; 
		5334: oled_colour = 16'b00001_000001_00001; 
		5335: oled_colour = 16'b00001_000001_00001; 
		5336: oled_colour = 16'b00001_000001_00001; 
		5337: oled_colour = 16'b00001_000001_00001; 
		5338: oled_colour = 16'b00001_000001_00001; 
		5339: oled_colour = 16'b00001_000001_00001; 
		5340: oled_colour = 16'b00001_000001_00001; 
		5341: oled_colour = 16'b00001_000001_00001; 
		5342: oled_colour = 16'b00001_000001_00001; 
		5343: oled_colour = 16'b00001_000001_00001; 
		5344: oled_colour = 16'b00001_000001_00001; 
		5345: oled_colour = 16'b00001_000001_00001; 
		5346: oled_colour = 16'b00001_000001_00001; 
		5347: oled_colour = 16'b00001_000001_00001; 
		5348: oled_colour = 16'b00001_000001_00001; 
		5349: oled_colour = 16'b00001_000001_00001; 
		5350: oled_colour = 16'b00001_000001_00001; 
		5351: oled_colour = 16'b00001_000001_00001; 
		5352: oled_colour = 16'b00001_000001_00001; 
		5353: oled_colour = 16'b00001_000001_00001; 
		5354: oled_colour = 16'b00001_000001_00001; 
		5355: oled_colour = 16'b00001_000001_00001; 
		5356: oled_colour = 16'b00001_000001_00001; 
		5357: oled_colour = 16'b00001_000001_00001; 
		5358: oled_colour = 16'b00001_000001_00001; 
		5359: oled_colour = 16'b00001_000001_00001; 
		5360: oled_colour = 16'b00001_000001_00001; 
		5361: oled_colour = 16'b00001_000001_00001; 
		5362: oled_colour = 16'b00001_000001_00001; 
		5363: oled_colour = 16'b00001_000001_00001; 
		5364: oled_colour = 16'b00001_000001_00001; 
		5365: oled_colour = 16'b00001_000001_00001; 
		5366: oled_colour = 16'b00001_000001_00001; 
		5367: oled_colour = 16'b00001_000001_00001; 
		5368: oled_colour = 16'b00001_000001_00001; 
		5369: oled_colour = 16'b00001_000001_00001; 
		5370: oled_colour = 16'b00001_000001_00001; 
		5371: oled_colour = 16'b00001_000001_00001; 
		5372: oled_colour = 16'b00001_000001_00001; 
		5373: oled_colour = 16'b00001_000001_00001; 
		5374: oled_colour = 16'b00001_000001_00001; 
		5375: oled_colour = 16'b00001_000001_00001; 
		5376: oled_colour = 16'b00001_000001_00001; 
		5377: oled_colour = 16'b00001_000001_00001; 
		5378: oled_colour = 16'b00001_000001_00001; 
		5379: oled_colour = 16'b00001_000001_00001; 
		5380: oled_colour = 16'b00001_000001_00001; 
		5381: oled_colour = 16'b00001_000001_00001; 
		5382: oled_colour = 16'b00001_000001_00001; 
		5383: oled_colour = 16'b00001_000001_00001; 
		5384: oled_colour = 16'b00001_000001_00001; 
		5385: oled_colour = 16'b00001_000001_00001; 
		5386: oled_colour = 16'b00001_000001_00001; 
		5387: oled_colour = 16'b00001_000001_00001; 
		5388: oled_colour = 16'b00001_000001_00001; 
		5389: oled_colour = 16'b00001_000001_00001; 
		5390: oled_colour = 16'b00001_000001_00001; 
		5391: oled_colour = 16'b00001_000001_00001; 
		5392: oled_colour = 16'b00001_000001_00001; 
		5393: oled_colour = 16'b00001_000001_00001; 
		5394: oled_colour = 16'b00001_000001_00001; 
		5395: oled_colour = 16'b00001_000001_00001; 
		5396: oled_colour = 16'b00001_000001_00001; 
		5397: oled_colour = 16'b00001_000001_00001; 
		5398: oled_colour = 16'b00001_000001_00001; 
		5399: oled_colour = 16'b00001_000001_00001; 
		5400: oled_colour = 16'b00001_000001_00001; 
		5401: oled_colour = 16'b00001_000001_00001; 
		5402: oled_colour = 16'b00001_000001_00001; 
		5403: oled_colour = 16'b00001_000001_00001; 
		5404: oled_colour = 16'b00001_000001_00001; 
		5405: oled_colour = 16'b00001_000001_00001; 
		5406: oled_colour = 16'b00001_000001_00001; 
		5407: oled_colour = 16'b00001_000001_00001; 
		5408: oled_colour = 16'b00001_000001_00001; 
		5409: oled_colour = 16'b00001_000001_00001; 
		5410: oled_colour = 16'b00001_000001_00001; 
		5411: oled_colour = 16'b00001_000001_00001; 
		5412: oled_colour = 16'b00001_000001_00001; 
		5413: oled_colour = 16'b00001_000001_00001; 
		5414: oled_colour = 16'b00001_000001_00001; 
		5415: oled_colour = 16'b00001_000001_00001; 
		5416: oled_colour = 16'b00001_000001_00001; 
		5417: oled_colour = 16'b00001_000001_00001; 
		5418: oled_colour = 16'b00001_000001_00001; 
		5419: oled_colour = 16'b00001_000001_00001; 
		5420: oled_colour = 16'b00001_000001_00001; 
		5421: oled_colour = 16'b00001_000001_00001; 
		5422: oled_colour = 16'b00001_000001_00001; 
		5423: oled_colour = 16'b00001_000001_00001; 
		5424: oled_colour = 16'b00001_000001_00001; 
		5425: oled_colour = 16'b00001_000001_00001; 
		5426: oled_colour = 16'b00001_000001_00001; 
		5427: oled_colour = 16'b00001_000001_00001; 
		5428: oled_colour = 16'b00001_000001_00001; 
		5429: oled_colour = 16'b00001_000001_00001; 
		5430: oled_colour = 16'b00001_000001_00001; 
		5431: oled_colour = 16'b00001_000001_00001; 
		5432: oled_colour = 16'b00001_000001_00001; 
		5433: oled_colour = 16'b00001_000001_00001; 
		5434: oled_colour = 16'b00001_000001_00001; 
		5435: oled_colour = 16'b00001_000001_00001; 
		5436: oled_colour = 16'b00001_000001_00001; 
		5437: oled_colour = 16'b00001_000001_00001; 
		5438: oled_colour = 16'b00001_000001_00001; 
		5439: oled_colour = 16'b00001_000001_00001; 
		5440: oled_colour = 16'b00001_000001_00001; 
		5441: oled_colour = 16'b00001_000001_00001; 
		5442: oled_colour = 16'b00001_000001_00001; 
		5443: oled_colour = 16'b00001_000001_00001; 
		5444: oled_colour = 16'b00001_000001_00001; 
		5445: oled_colour = 16'b00001_000001_00001; 
		5446: oled_colour = 16'b00001_000001_00001; 
		5447: oled_colour = 16'b00001_000001_00001; 
		5448: oled_colour = 16'b00001_000001_00001; 
		5449: oled_colour = 16'b00001_000001_00001; 
		5450: oled_colour = 16'b00001_000001_00001; 
		5451: oled_colour = 16'b00001_000001_00001; 
		5452: oled_colour = 16'b00001_000001_00001; 
		5453: oled_colour = 16'b00001_000001_00001; 
		5454: oled_colour = 16'b00001_000001_00001; 
		5455: oled_colour = 16'b00001_000001_00001; 
		5456: oled_colour = 16'b00001_000001_00001; 
		5457: oled_colour = 16'b00001_000001_00001; 
		5458: oled_colour = 16'b00001_000001_00001; 
		5459: oled_colour = 16'b00001_000001_00001; 
		5460: oled_colour = 16'b00001_000001_00001; 
		5461: oled_colour = 16'b00001_000001_00001; 
		5462: oled_colour = 16'b00001_000001_00001; 
		5463: oled_colour = 16'b00001_000001_00001; 
		5464: oled_colour = 16'b00001_000001_00001; 
		5465: oled_colour = 16'b00001_000001_00001; 
		5466: oled_colour = 16'b00001_000001_00001; 
		5467: oled_colour = 16'b00001_000001_00001; 
		5468: oled_colour = 16'b00001_000001_00001; 
		5469: oled_colour = 16'b00001_000001_00001; 
		5470: oled_colour = 16'b00001_000001_00001; 
		5471: oled_colour = 16'b00001_000001_00001; 
		5472: oled_colour = 16'b00001_000001_00001; 
		5473: oled_colour = 16'b00001_000001_00001; 
		5474: oled_colour = 16'b00001_000001_00001; 
		5475: oled_colour = 16'b00001_000001_00001; 
		5476: oled_colour = 16'b00001_000001_00001; 
		5477: oled_colour = 16'b00001_000001_00001; 
		5478: oled_colour = 16'b00001_000001_00001; 
		5479: oled_colour = 16'b00001_000001_00001; 
		5480: oled_colour = 16'b00001_000001_00001; 
		5481: oled_colour = 16'b00001_000001_00001; 
		5482: oled_colour = 16'b00001_000001_00001; 
		5483: oled_colour = 16'b00001_000001_00001; 
		5484: oled_colour = 16'b00001_000001_00001; 
		5485: oled_colour = 16'b00001_000001_00001; 
		5486: oled_colour = 16'b00001_000001_00001; 
		5487: oled_colour = 16'b00001_000001_00001; 
		5488: oled_colour = 16'b00001_000001_00001; 
		5489: oled_colour = 16'b00001_000001_00001; 
		5490: oled_colour = 16'b00001_000001_00001; 
		5491: oled_colour = 16'b00001_000001_00001; 
		5492: oled_colour = 16'b00001_000001_00001; 
		5493: oled_colour = 16'b00001_000001_00001; 
		5494: oled_colour = 16'b00001_000001_00001; 
		5495: oled_colour = 16'b00001_000001_00001; 
		5496: oled_colour = 16'b00001_000001_00001; 
		5497: oled_colour = 16'b00001_000001_00001; 
		5498: oled_colour = 16'b00001_000001_00001; 
		5499: oled_colour = 16'b00001_000001_00001; 
		5500: oled_colour = 16'b00001_000001_00001; 
		5501: oled_colour = 16'b00001_000001_00001; 
		5502: oled_colour = 16'b00001_000001_00001; 
		5503: oled_colour = 16'b00001_000001_00001; 
		5504: oled_colour = 16'b00001_000001_00001; 
		5505: oled_colour = 16'b00001_000001_00001; 
		5506: oled_colour = 16'b00001_000001_00001; 
		5507: oled_colour = 16'b00001_000001_00001; 
		5508: oled_colour = 16'b00001_000001_00001; 
		5509: oled_colour = 16'b00001_000001_00001; 
		5510: oled_colour = 16'b00001_000001_00001; 
		5511: oled_colour = 16'b00001_000001_00001; 
		5512: oled_colour = 16'b00001_000001_00001; 
		5513: oled_colour = 16'b00001_000001_00001; 
		5514: oled_colour = 16'b00001_000001_00001; 
		5515: oled_colour = 16'b00001_000001_00001; 
		5516: oled_colour = 16'b00001_000001_00001; 
		5517: oled_colour = 16'b00001_000001_00001; 
		5518: oled_colour = 16'b00001_000001_00001; 
		5519: oled_colour = 16'b00001_000001_00001; 
		5520: oled_colour = 16'b00001_000001_00001; 
		5521: oled_colour = 16'b00001_000001_00001; 
		5522: oled_colour = 16'b00001_000001_00001; 
		5523: oled_colour = 16'b00001_000001_00001; 
		5524: oled_colour = 16'b00001_000001_00001; 
		5525: oled_colour = 16'b00001_000001_00001; 
		5526: oled_colour = 16'b00001_000001_00001; 
		5527: oled_colour = 16'b00001_000001_00001; 
		5528: oled_colour = 16'b00001_000001_00001; 
		5529: oled_colour = 16'b00001_000001_00001; 
		5530: oled_colour = 16'b00001_000001_00001; 
		5531: oled_colour = 16'b00001_000001_00001; 
		5532: oled_colour = 16'b00001_000001_00001; 
		5533: oled_colour = 16'b00001_000001_00001; 
		5534: oled_colour = 16'b00001_000001_00001; 
		5535: oled_colour = 16'b00001_000001_00001; 
		5536: oled_colour = 16'b00001_000001_00001; 
		5537: oled_colour = 16'b00001_000001_00001; 
		5538: oled_colour = 16'b00001_000001_00001; 
		5539: oled_colour = 16'b00001_000001_00001; 
		5540: oled_colour = 16'b00001_000001_00001; 
		5541: oled_colour = 16'b00001_000001_00001; 
		5542: oled_colour = 16'b00001_000001_00001; 
		5543: oled_colour = 16'b00001_000001_00001; 
		5544: oled_colour = 16'b00001_000001_00001; 
		5545: oled_colour = 16'b00001_000001_00001; 
		5546: oled_colour = 16'b00001_000001_00001; 
		5547: oled_colour = 16'b00001_000001_00001; 
		5548: oled_colour = 16'b00001_000001_00001; 
		5549: oled_colour = 16'b00001_000001_00001; 
		5550: oled_colour = 16'b00001_000001_00001; 
		5551: oled_colour = 16'b00001_000001_00001; 
		5552: oled_colour = 16'b00001_000001_00001; 
		5553: oled_colour = 16'b00001_000001_00001; 
		5554: oled_colour = 16'b00001_000001_00001; 
		5555: oled_colour = 16'b00001_000001_00001; 
		5556: oled_colour = 16'b00001_000001_00001; 
		5557: oled_colour = 16'b00001_000001_00001; 
		5558: oled_colour = 16'b00001_000001_00001; 
		5559: oled_colour = 16'b00001_000001_00001; 
		5560: oled_colour = 16'b00001_000001_00001; 
		5561: oled_colour = 16'b00001_000001_00001; 
		5562: oled_colour = 16'b00001_000001_00001; 
		5563: oled_colour = 16'b00001_000001_00001; 
		5564: oled_colour = 16'b00001_000001_00001; 
		5565: oled_colour = 16'b00001_000001_00001; 
		5566: oled_colour = 16'b00001_000001_00001; 
		5567: oled_colour = 16'b00001_000001_00001; 
		5568: oled_colour = 16'b00001_000001_00001; 
		5569: oled_colour = 16'b00001_000001_00001; 
		5570: oled_colour = 16'b00001_000001_00001; 
		5571: oled_colour = 16'b00001_000001_00001; 
		5572: oled_colour = 16'b00001_000001_00001; 
		5573: oled_colour = 16'b00001_000001_00001; 
		5574: oled_colour = 16'b00001_000001_00001; 
		5575: oled_colour = 16'b00001_000001_00001; 
		5576: oled_colour = 16'b00001_000001_00001; 
		5577: oled_colour = 16'b00001_000001_00001; 
		5578: oled_colour = 16'b00001_000001_00001; 
		5579: oled_colour = 16'b00001_000001_00001; 
		5580: oled_colour = 16'b00001_000001_00001; 
		5581: oled_colour = 16'b00001_000001_00001; 
		5582: oled_colour = 16'b00001_000001_00001; 
		5583: oled_colour = 16'b00001_000001_00001; 
		5584: oled_colour = 16'b00001_000001_00001; 
		5585: oled_colour = 16'b00001_000001_00001; 
		5586: oled_colour = 16'b00001_000001_00001; 
		5587: oled_colour = 16'b00001_000001_00001; 
		5588: oled_colour = 16'b00001_000001_00001; 
		5589: oled_colour = 16'b00001_000001_00001; 
		5590: oled_colour = 16'b00001_000001_00001; 
		5591: oled_colour = 16'b00001_000001_00001; 
		5592: oled_colour = 16'b00001_000001_00001; 
		5593: oled_colour = 16'b00001_000001_00001; 
		5594: oled_colour = 16'b00001_000001_00001; 
		5595: oled_colour = 16'b00001_000001_00001; 
		5596: oled_colour = 16'b00001_000001_00001; 
		5597: oled_colour = 16'b00001_000001_00001; 
		5598: oled_colour = 16'b00001_000001_00001; 
		5599: oled_colour = 16'b00001_000001_00001; 
		5600: oled_colour = 16'b00001_000001_00001; 
		5601: oled_colour = 16'b00001_000001_00001; 
		5602: oled_colour = 16'b00001_000001_00001; 
		5603: oled_colour = 16'b00001_000001_00001; 
		5604: oled_colour = 16'b00001_000001_00001; 
		5605: oled_colour = 16'b00001_000001_00001; 
		5606: oled_colour = 16'b00001_000001_00001; 
		5607: oled_colour = 16'b00001_000001_00001; 
		5608: oled_colour = 16'b00001_000001_00001; 
		5609: oled_colour = 16'b00001_000001_00001; 
		5610: oled_colour = 16'b00001_000001_00001; 
		5611: oled_colour = 16'b00001_000001_00001; 
		5612: oled_colour = 16'b00001_000001_00001; 
		5613: oled_colour = 16'b00001_000001_00001; 
		5614: oled_colour = 16'b00001_000001_00001; 
		5615: oled_colour = 16'b00001_000001_00001; 
		5616: oled_colour = 16'b00001_000001_00001; 
		5617: oled_colour = 16'b00001_000001_00001; 
		5618: oled_colour = 16'b00001_000001_00001; 
		5619: oled_colour = 16'b00001_000001_00001; 
		5620: oled_colour = 16'b00001_000001_00001; 
		5621: oled_colour = 16'b00001_000001_00001; 
		5622: oled_colour = 16'b00001_000001_00001; 
		5623: oled_colour = 16'b00001_000001_00001; 
		5624: oled_colour = 16'b00001_000001_00001; 
		5625: oled_colour = 16'b00001_000001_00001; 
		5626: oled_colour = 16'b00001_000001_00001; 
		5627: oled_colour = 16'b00001_000001_00001; 
		5628: oled_colour = 16'b00001_000001_00001; 
		5629: oled_colour = 16'b00001_000001_00001; 
		5630: oled_colour = 16'b00001_000001_00001; 
		5631: oled_colour = 16'b00001_000001_00001; 
		5632: oled_colour = 16'b00001_000001_00001; 
		5633: oled_colour = 16'b00001_000001_00001; 
		5634: oled_colour = 16'b00001_000001_00001; 
		5635: oled_colour = 16'b00001_000001_00001; 
		5636: oled_colour = 16'b00001_000001_00001; 
		5637: oled_colour = 16'b00001_000001_00001; 
		5638: oled_colour = 16'b00001_000001_00001; 
		5639: oled_colour = 16'b00001_000001_00001; 
		5640: oled_colour = 16'b00001_000001_00001; 
		5641: oled_colour = 16'b00001_000001_00001; 
		5642: oled_colour = 16'b00001_000001_00001; 
		5643: oled_colour = 16'b00001_000001_00001; 
		5644: oled_colour = 16'b00001_000001_00001; 
		5645: oled_colour = 16'b00001_000001_00001; 
		5646: oled_colour = 16'b00001_000001_00001; 
		5647: oled_colour = 16'b00001_000001_00001; 
		5648: oled_colour = 16'b00001_000001_00001; 
		5649: oled_colour = 16'b00001_000001_00001; 
		5650: oled_colour = 16'b00001_000001_00001; 
		5651: oled_colour = 16'b00001_000001_00001; 
		5652: oled_colour = 16'b00001_000001_00001; 
		5653: oled_colour = 16'b00001_000001_00001; 
		5654: oled_colour = 16'b00001_000001_00001; 
		5655: oled_colour = 16'b00001_000001_00001; 
		5656: oled_colour = 16'b00001_000001_00001; 
		5657: oled_colour = 16'b00001_000001_00001; 
		5658: oled_colour = 16'b00001_000001_00001; 
		5659: oled_colour = 16'b00001_000001_00001; 
		5660: oled_colour = 16'b00001_000001_00001; 
		5661: oled_colour = 16'b00001_000001_00001; 
		5662: oled_colour = 16'b00001_000001_00001; 
		5663: oled_colour = 16'b00001_000001_00001; 
		5664: oled_colour = 16'b00001_000001_00001; 
		5665: oled_colour = 16'b00001_000001_00001; 
		5666: oled_colour = 16'b00001_000001_00001; 
		5667: oled_colour = 16'b00001_000001_00001; 
		5668: oled_colour = 16'b00001_000001_00001; 
		5669: oled_colour = 16'b00001_000001_00001; 
		5670: oled_colour = 16'b00001_000001_00001; 
		5671: oled_colour = 16'b00001_000001_00001; 
		5672: oled_colour = 16'b00001_000001_00001; 
		5673: oled_colour = 16'b00001_000001_00001; 
		5674: oled_colour = 16'b00001_000001_00001; 
		5675: oled_colour = 16'b00001_000001_00001; 
		5676: oled_colour = 16'b00001_000001_00001; 
		5677: oled_colour = 16'b00001_000001_00001; 
		5678: oled_colour = 16'b00001_000001_00001; 
		5679: oled_colour = 16'b00001_000001_00001; 
		5680: oled_colour = 16'b00001_000001_00001; 
		5681: oled_colour = 16'b00001_000001_00001; 
		5682: oled_colour = 16'b00001_000001_00001; 
		5683: oled_colour = 16'b00001_000001_00001; 
		5684: oled_colour = 16'b00001_000001_00001; 
		5685: oled_colour = 16'b00001_000001_00001; 
		5686: oled_colour = 16'b00001_000001_00001; 
		5687: oled_colour = 16'b00001_000001_00001; 
		5688: oled_colour = 16'b00001_000001_00001; 
		5689: oled_colour = 16'b00001_000001_00001; 
		5690: oled_colour = 16'b00001_000001_00001; 
		5691: oled_colour = 16'b00001_000001_00001; 
		5692: oled_colour = 16'b00001_000001_00001; 
		5693: oled_colour = 16'b00001_000001_00001; 
		5694: oled_colour = 16'b00001_000001_00001; 
		5695: oled_colour = 16'b00001_000001_00001; 
		5696: oled_colour = 16'b00001_000001_00001; 
		5697: oled_colour = 16'b00001_000001_00001; 
		5698: oled_colour = 16'b00001_000001_00001; 
		5699: oled_colour = 16'b00001_000001_00001; 
		5700: oled_colour = 16'b00001_000001_00001; 
		5701: oled_colour = 16'b00001_000001_00001; 
		5702: oled_colour = 16'b00001_000001_00001; 
		5703: oled_colour = 16'b00001_000001_00001; 
		5704: oled_colour = 16'b00001_000001_00001; 
		5705: oled_colour = 16'b00001_000001_00001; 
		5706: oled_colour = 16'b00001_000001_00001; 
		5707: oled_colour = 16'b00001_000001_00001; 
		5708: oled_colour = 16'b00001_000001_00001; 
		5709: oled_colour = 16'b00001_000001_00001; 
		5710: oled_colour = 16'b00001_000001_00001; 
		5711: oled_colour = 16'b00001_000001_00001; 
		5712: oled_colour = 16'b00001_000001_00001; 
		5713: oled_colour = 16'b00001_000001_00001; 
		5714: oled_colour = 16'b00001_000001_00001; 
		5715: oled_colour = 16'b00001_000001_00001; 
		5716: oled_colour = 16'b00001_000001_00001; 
		5717: oled_colour = 16'b00001_000001_00001; 
		5718: oled_colour = 16'b00001_000001_00001; 
		5719: oled_colour = 16'b00001_000001_00001; 
		5720: oled_colour = 16'b00001_000001_00001; 
		5721: oled_colour = 16'b00001_000001_00001; 
		5722: oled_colour = 16'b00001_000001_00001; 
		5723: oled_colour = 16'b00001_000001_00001; 
		5724: oled_colour = 16'b00001_000001_00001; 
		5725: oled_colour = 16'b00001_000001_00001; 
		5726: oled_colour = 16'b00001_000001_00001; 
		5727: oled_colour = 16'b00001_000001_00001; 
		5728: oled_colour = 16'b00001_000001_00001; 
		5729: oled_colour = 16'b00001_000001_00001; 
		5730: oled_colour = 16'b00001_000001_00001; 
		5731: oled_colour = 16'b00001_000001_00001; 
		5732: oled_colour = 16'b00001_000001_00001; 
		5733: oled_colour = 16'b00001_000001_00001; 
		5734: oled_colour = 16'b00001_000001_00001; 
		5735: oled_colour = 16'b00001_000001_00001; 
		5736: oled_colour = 16'b00001_000001_00001; 
		5737: oled_colour = 16'b00001_000001_00001; 
		5738: oled_colour = 16'b00001_000001_00001; 
		5739: oled_colour = 16'b00001_000001_00001; 
		5740: oled_colour = 16'b00001_000001_00001; 
		5741: oled_colour = 16'b00001_000001_00001; 
		5742: oled_colour = 16'b00001_000001_00001; 
		5743: oled_colour = 16'b00001_000001_00001; 
		5744: oled_colour = 16'b00001_000001_00001; 
		5745: oled_colour = 16'b00001_000001_00001; 
		5746: oled_colour = 16'b00001_000001_00001; 
		5747: oled_colour = 16'b00001_000001_00001; 
		5748: oled_colour = 16'b00001_000001_00001; 
		5749: oled_colour = 16'b00001_000001_00001; 
		5750: oled_colour = 16'b00001_000001_00001; 
		5751: oled_colour = 16'b00001_000001_00001; 
		5752: oled_colour = 16'b00001_000001_00001; 
		5753: oled_colour = 16'b00001_000001_00001; 
		5754: oled_colour = 16'b00001_000001_00001; 
		5755: oled_colour = 16'b00001_000001_00001; 
		5756: oled_colour = 16'b00001_000001_00001; 
		5757: oled_colour = 16'b00001_000001_00001; 
		5758: oled_colour = 16'b00001_000001_00001; 
		5759: oled_colour = 16'b00001_000001_00001; 
		5760: oled_colour = 16'b00001_000001_00001; 
		5761: oled_colour = 16'b00001_000001_00001; 
		5762: oled_colour = 16'b00001_000001_00001; 
		5763: oled_colour = 16'b00001_000001_00001; 
		5764: oled_colour = 16'b00001_000001_00001; 
		5765: oled_colour = 16'b00001_000001_00001; 
		5766: oled_colour = 16'b00001_000001_00001; 
		5767: oled_colour = 16'b00001_000001_00001; 
		5768: oled_colour = 16'b00001_000001_00001; 
		5769: oled_colour = 16'b00001_000001_00001; 
		5770: oled_colour = 16'b00001_000001_00001; 
		5771: oled_colour = 16'b00001_000001_00001; 
		5772: oled_colour = 16'b00001_000001_00001; 
		5773: oled_colour = 16'b00001_000001_00001; 
		5774: oled_colour = 16'b00001_000001_00001; 
		5775: oled_colour = 16'b00001_000001_00001; 
		5776: oled_colour = 16'b00001_000001_00001; 
		5777: oled_colour = 16'b00001_000001_00001; 
		5778: oled_colour = 16'b00001_000001_00001; 
		5779: oled_colour = 16'b00001_000001_00001; 
		5780: oled_colour = 16'b00001_000001_00001; 
		5781: oled_colour = 16'b00001_000001_00001; 
		5782: oled_colour = 16'b00001_000001_00001; 
		5783: oled_colour = 16'b00001_000001_00001; 
		5784: oled_colour = 16'b00001_000001_00001; 
		5785: oled_colour = 16'b00001_000001_00001; 
		5786: oled_colour = 16'b00001_000001_00001; 
		5787: oled_colour = 16'b00001_000001_00001; 
		5788: oled_colour = 16'b00001_000001_00001; 
		5789: oled_colour = 16'b00001_000001_00001; 
		5790: oled_colour = 16'b00001_000001_00001; 
		5791: oled_colour = 16'b00001_000001_00001; 
		5792: oled_colour = 16'b00001_000001_00001; 
		5793: oled_colour = 16'b00001_000001_00001; 
		5794: oled_colour = 16'b00001_000001_00001; 
		5795: oled_colour = 16'b00001_000001_00001; 
		5796: oled_colour = 16'b00001_000001_00001; 
		5797: oled_colour = 16'b00001_000001_00001; 
		5798: oled_colour = 16'b00001_000001_00001; 
		5799: oled_colour = 16'b00001_000001_00001; 
		5800: oled_colour = 16'b00001_000001_00001; 
		5801: oled_colour = 16'b00001_000001_00001; 
		5802: oled_colour = 16'b00001_000001_00001; 
		5803: oled_colour = 16'b00001_000001_00001; 
		5804: oled_colour = 16'b00001_000001_00001; 
		5805: oled_colour = 16'b00001_000001_00001; 
		5806: oled_colour = 16'b00001_000001_00001; 
		5807: oled_colour = 16'b00001_000001_00001; 
		5808: oled_colour = 16'b00001_000001_00001; 
		5809: oled_colour = 16'b00001_000001_00001; 
		5810: oled_colour = 16'b00001_000001_00001; 
		5811: oled_colour = 16'b00001_000001_00001; 
		5812: oled_colour = 16'b00001_000001_00001; 
		5813: oled_colour = 16'b00001_000001_00001; 
		5814: oled_colour = 16'b00001_000001_00001; 
		5815: oled_colour = 16'b00001_000001_00001; 
		5816: oled_colour = 16'b00001_000001_00001; 
		5817: oled_colour = 16'b00001_000001_00001; 
		5818: oled_colour = 16'b00001_000001_00001; 
		5819: oled_colour = 16'b00001_000001_00001; 
		5820: oled_colour = 16'b00001_000001_00001; 
		5821: oled_colour = 16'b00001_000001_00001; 
		5822: oled_colour = 16'b00001_000001_00001; 
		5823: oled_colour = 16'b00001_000001_00001; 
		5824: oled_colour = 16'b00001_000001_00001; 
		5825: oled_colour = 16'b00001_000001_00001; 
		5826: oled_colour = 16'b00001_000001_00001; 
		5827: oled_colour = 16'b00001_000001_00001; 
		5828: oled_colour = 16'b00001_000001_00001; 
		5829: oled_colour = 16'b00001_000001_00001; 
		5830: oled_colour = 16'b00001_000001_00001; 
		5831: oled_colour = 16'b00001_000001_00001; 
		5832: oled_colour = 16'b00001_000001_00001; 
		5833: oled_colour = 16'b00001_000001_00001; 
		5834: oled_colour = 16'b00001_000001_00001; 
		5835: oled_colour = 16'b00001_000001_00001; 
		5836: oled_colour = 16'b00001_000001_00001; 
		5837: oled_colour = 16'b00001_000001_00001; 
		5838: oled_colour = 16'b00001_000001_00001; 
		5839: oled_colour = 16'b00001_000001_00001; 
		5840: oled_colour = 16'b00001_000001_00001; 
		5841: oled_colour = 16'b00001_000001_00001; 
		5842: oled_colour = 16'b00001_000001_00001; 
		5843: oled_colour = 16'b00001_000001_00001; 
		5844: oled_colour = 16'b00001_000001_00001; 
		5845: oled_colour = 16'b00001_000001_00001; 
		5846: oled_colour = 16'b00001_000001_00001; 
		5847: oled_colour = 16'b00001_000001_00001; 
		5848: oled_colour = 16'b00001_000001_00001; 
		5849: oled_colour = 16'b00001_000001_00001; 
		5850: oled_colour = 16'b00001_000001_00001; 
		5851: oled_colour = 16'b00001_000001_00001; 
		5852: oled_colour = 16'b00001_000001_00001; 
		5853: oled_colour = 16'b00001_000001_00001; 
		5854: oled_colour = 16'b00001_000001_00001; 
		5855: oled_colour = 16'b00001_000001_00001; 
		5856: oled_colour = 16'b00001_000001_00001; 
		5857: oled_colour = 16'b00001_000001_00001; 
		5858: oled_colour = 16'b00001_000001_00001; 
		5859: oled_colour = 16'b00001_000001_00001; 
		5860: oled_colour = 16'b00001_000001_00001; 
		5861: oled_colour = 16'b00001_000001_00001; 
		5862: oled_colour = 16'b00001_000001_00001; 
		5863: oled_colour = 16'b00001_000001_00001; 
		5864: oled_colour = 16'b00001_000001_00001; 
		5865: oled_colour = 16'b00001_000001_00001; 
		5866: oled_colour = 16'b00001_000001_00001; 
		5867: oled_colour = 16'b00001_000001_00001; 
		5868: oled_colour = 16'b00001_000001_00001; 
		5869: oled_colour = 16'b00001_000001_00001; 
		5870: oled_colour = 16'b00001_000001_00001; 
		5871: oled_colour = 16'b00001_000001_00001; 
		5872: oled_colour = 16'b00001_000001_00001; 
		5873: oled_colour = 16'b00001_000001_00001; 
		5874: oled_colour = 16'b00001_000001_00001; 
		5875: oled_colour = 16'b00001_000001_00001; 
		5876: oled_colour = 16'b00001_000001_00001; 
		5877: oled_colour = 16'b00001_000001_00001; 
		5878: oled_colour = 16'b00001_000001_00001; 
		5879: oled_colour = 16'b00001_000001_00001; 
		5880: oled_colour = 16'b00001_000001_00001; 
		5881: oled_colour = 16'b00001_000001_00001; 
		5882: oled_colour = 16'b00001_000001_00001; 
		5883: oled_colour = 16'b00001_000001_00001; 
		5884: oled_colour = 16'b00001_000001_00001; 
		5885: oled_colour = 16'b00001_000001_00001; 
		5886: oled_colour = 16'b00001_000001_00001; 
		5887: oled_colour = 16'b00001_000001_00001; 
		5888: oled_colour = 16'b00001_000001_00001; 
		5889: oled_colour = 16'b00001_000001_00001; 
		5890: oled_colour = 16'b00001_000001_00001; 
		5891: oled_colour = 16'b00001_000001_00001; 
		5892: oled_colour = 16'b00001_000001_00001; 
		5893: oled_colour = 16'b00001_000001_00001; 
		5894: oled_colour = 16'b00001_000001_00001; 
		5895: oled_colour = 16'b00001_000001_00001; 
		5896: oled_colour = 16'b00001_000001_00001; 
		5897: oled_colour = 16'b00001_000001_00001; 
		5898: oled_colour = 16'b00001_000001_00001; 
		5899: oled_colour = 16'b00001_000001_00001; 
		5900: oled_colour = 16'b00001_000001_00001; 
		5901: oled_colour = 16'b00001_000001_00001; 
		5902: oled_colour = 16'b00001_000001_00001; 
		5903: oled_colour = 16'b00001_000001_00001; 
		5904: oled_colour = 16'b00001_000001_00001; 
		5905: oled_colour = 16'b00001_000001_00001; 
		5906: oled_colour = 16'b00001_000001_00001; 
		5907: oled_colour = 16'b00001_000001_00001; 
		5908: oled_colour = 16'b00001_000001_00001; 
		5909: oled_colour = 16'b00001_000001_00001; 
		5910: oled_colour = 16'b00001_000001_00001; 
		5911: oled_colour = 16'b00001_000001_00001; 
		5912: oled_colour = 16'b00001_000001_00001; 
		5913: oled_colour = 16'b00001_000001_00001; 
		5914: oled_colour = 16'b00001_000001_00001; 
		5915: oled_colour = 16'b00001_000001_00001; 
		5916: oled_colour = 16'b00001_000001_00001; 
		5917: oled_colour = 16'b00001_000001_00001; 
		5918: oled_colour = 16'b00001_000001_00001; 
		5919: oled_colour = 16'b00001_000001_00001; 
		5920: oled_colour = 16'b00001_000001_00001; 
		5921: oled_colour = 16'b00001_000001_00001; 
		5922: oled_colour = 16'b00001_000001_00001; 
		5923: oled_colour = 16'b00001_000001_00001; 
		5924: oled_colour = 16'b00001_000001_00001; 
		5925: oled_colour = 16'b00001_000001_00001; 
		5926: oled_colour = 16'b00001_000001_00001; 
		5927: oled_colour = 16'b00001_000001_00001; 
		5928: oled_colour = 16'b00001_000001_00001; 
		5929: oled_colour = 16'b00001_000001_00001; 
		5930: oled_colour = 16'b00001_000001_00001; 
		5931: oled_colour = 16'b00001_000001_00001; 
		5932: oled_colour = 16'b00001_000001_00001; 
		5933: oled_colour = 16'b00001_000001_00001; 
		5934: oled_colour = 16'b00001_000001_00001; 
		5935: oled_colour = 16'b00001_000001_00001; 
		5936: oled_colour = 16'b00001_000001_00001; 
		5937: oled_colour = 16'b00001_000001_00001; 
		5938: oled_colour = 16'b00001_000001_00001; 
		5939: oled_colour = 16'b00001_000001_00001; 
		5940: oled_colour = 16'b00001_000001_00001; 
		5941: oled_colour = 16'b00001_000001_00001; 
		5942: oled_colour = 16'b00001_000001_00001; 
		5943: oled_colour = 16'b00001_000001_00001; 
		5944: oled_colour = 16'b00001_000001_00001; 
		5945: oled_colour = 16'b00001_000001_00001; 
		5946: oled_colour = 16'b00001_000001_00001; 
		5947: oled_colour = 16'b00001_000001_00001; 
		5948: oled_colour = 16'b00001_000001_00001; 
		5949: oled_colour = 16'b00001_000001_00001; 
		5950: oled_colour = 16'b00001_000001_00001; 
		5951: oled_colour = 16'b00001_000001_00001; 
		5952: oled_colour = 16'b00001_000001_00001; 
		5953: oled_colour = 16'b00001_000001_00001; 
		5954: oled_colour = 16'b00001_000001_00001; 
		5955: oled_colour = 16'b00001_000001_00001; 
		5956: oled_colour = 16'b00001_000001_00001; 
		5957: oled_colour = 16'b00001_000001_00001; 
		5958: oled_colour = 16'b00001_000001_00001; 
		5959: oled_colour = 16'b00001_000001_00001; 
		5960: oled_colour = 16'b00001_000001_00001; 
		5961: oled_colour = 16'b00001_000001_00001; 
		5962: oled_colour = 16'b00001_000001_00001; 
		5963: oled_colour = 16'b00001_000001_00001; 
		5964: oled_colour = 16'b00001_000001_00001; 
		5965: oled_colour = 16'b00001_000001_00001; 
		5966: oled_colour = 16'b00001_000001_00001; 
		5967: oled_colour = 16'b00001_000001_00001; 
		5968: oled_colour = 16'b00001_000001_00001; 
		5969: oled_colour = 16'b00001_000001_00001; 
		5970: oled_colour = 16'b00001_000001_00001; 
		5971: oled_colour = 16'b00001_000001_00001; 
		5972: oled_colour = 16'b00001_000001_00001; 
		5973: oled_colour = 16'b00001_000001_00001; 
		5974: oled_colour = 16'b00001_000001_00001; 
		5975: oled_colour = 16'b00001_000001_00001; 
		5976: oled_colour = 16'b00001_000001_00001; 
		5977: oled_colour = 16'b00001_000001_00001; 
		5978: oled_colour = 16'b00001_000001_00001; 
		5979: oled_colour = 16'b00001_000001_00001; 
		5980: oled_colour = 16'b00001_000001_00001; 
		5981: oled_colour = 16'b00001_000001_00001; 
		5982: oled_colour = 16'b00001_000001_00001; 
		5983: oled_colour = 16'b00001_000001_00001; 
		5984: oled_colour = 16'b00001_000001_00001; 
		5985: oled_colour = 16'b00001_000001_00001; 
		5986: oled_colour = 16'b00001_000001_00001; 
		5987: oled_colour = 16'b00001_000001_00001; 
		5988: oled_colour = 16'b00001_000001_00001; 
		5989: oled_colour = 16'b00001_000001_00001; 
		5990: oled_colour = 16'b00001_000001_00001; 
		5991: oled_colour = 16'b00001_000001_00001; 
		5992: oled_colour = 16'b00001_000001_00001; 
		5993: oled_colour = 16'b00001_000001_00001; 
		5994: oled_colour = 16'b00001_000001_00001; 
		5995: oled_colour = 16'b00001_000001_00001; 
		5996: oled_colour = 16'b00001_000001_00001; 
		5997: oled_colour = 16'b00001_000001_00001; 
		5998: oled_colour = 16'b00001_000001_00001; 
		5999: oled_colour = 16'b00001_000001_00001; 
		6000: oled_colour = 16'b00001_000001_00001; 
		6001: oled_colour = 16'b00001_000001_00001; 
		6002: oled_colour = 16'b00001_000001_00001; 
		6003: oled_colour = 16'b00001_000001_00001; 
		6004: oled_colour = 16'b00001_000001_00001; 
		6005: oled_colour = 16'b00001_000001_00001; 
		6006: oled_colour = 16'b00001_000001_00001; 
		6007: oled_colour = 16'b00001_000001_00001; 
		6008: oled_colour = 16'b00001_000001_00001; 
		6009: oled_colour = 16'b00001_000001_00001; 
		6010: oled_colour = 16'b00001_000001_00001; 
		6011: oled_colour = 16'b00001_000001_00001; 
		6012: oled_colour = 16'b00001_000001_00001; 
		6013: oled_colour = 16'b00001_000001_00001; 
		6014: oled_colour = 16'b00001_000001_00001; 
		6015: oled_colour = 16'b00001_000001_00001; 
		6016: oled_colour = 16'b00001_000001_00001; 
		6017: oled_colour = 16'b00001_000001_00001; 
		6018: oled_colour = 16'b00001_000001_00001; 
		6019: oled_colour = 16'b00001_000001_00001; 
		6020: oled_colour = 16'b00001_000001_00001; 
		6021: oled_colour = 16'b00001_000001_00001; 
		6022: oled_colour = 16'b00001_000001_00001; 
		6023: oled_colour = 16'b00001_000001_00001; 
		6024: oled_colour = 16'b00001_000001_00001; 
		6025: oled_colour = 16'b00001_000001_00001; 
		6026: oled_colour = 16'b00001_000001_00001; 
		6027: oled_colour = 16'b00001_000001_00001; 
		6028: oled_colour = 16'b00001_000001_00001; 
		6029: oled_colour = 16'b00001_000001_00001; 
		6030: oled_colour = 16'b00001_000001_00001; 
		6031: oled_colour = 16'b00001_000001_00001; 
		6032: oled_colour = 16'b00001_000001_00001; 
		6033: oled_colour = 16'b00001_000001_00001; 
		6034: oled_colour = 16'b00001_000001_00001; 
		6035: oled_colour = 16'b00001_000001_00001; 
		6036: oled_colour = 16'b00001_000001_00001; 
		6037: oled_colour = 16'b00001_000001_00001; 
		6038: oled_colour = 16'b00001_000001_00001; 
		6039: oled_colour = 16'b00001_000001_00001; 
		6040: oled_colour = 16'b00001_000001_00001; 
		6041: oled_colour = 16'b00001_000001_00001; 
		6042: oled_colour = 16'b00001_000001_00001; 
		6043: oled_colour = 16'b00001_000001_00001; 
		6044: oled_colour = 16'b00001_000001_00001; 
		6045: oled_colour = 16'b00001_000001_00001; 
		6046: oled_colour = 16'b00001_000001_00001; 
		6047: oled_colour = 16'b00001_000001_00001; 
		6048: oled_colour = 16'b00001_000001_00001; 
		6049: oled_colour = 16'b00001_000001_00001; 
		6050: oled_colour = 16'b00001_000001_00001; 
		6051: oled_colour = 16'b00001_000001_00001; 
		6052: oled_colour = 16'b00001_000001_00001; 
		6053: oled_colour = 16'b00001_000001_00001; 
		6054: oled_colour = 16'b00001_000001_00001; 
		6055: oled_colour = 16'b00001_000001_00001; 
		6056: oled_colour = 16'b00001_000001_00001; 
		6057: oled_colour = 16'b00001_000001_00001; 
		6058: oled_colour = 16'b00001_000001_00001; 
		6059: oled_colour = 16'b00001_000001_00001; 
		6060: oled_colour = 16'b00001_000001_00001; 
		6061: oled_colour = 16'b00001_000001_00001; 
		6062: oled_colour = 16'b00001_000001_00001; 
		6063: oled_colour = 16'b00001_000001_00001; 
		6064: oled_colour = 16'b00001_000001_00001; 
		6065: oled_colour = 16'b00001_000001_00001; 
		6066: oled_colour = 16'b00001_000001_00001; 
		6067: oled_colour = 16'b00001_000001_00001; 
		6068: oled_colour = 16'b00001_000001_00001; 
		6069: oled_colour = 16'b00001_000001_00001; 
		6070: oled_colour = 16'b00001_000001_00001; 
		6071: oled_colour = 16'b00001_000001_00001; 
		6072: oled_colour = 16'b00001_000001_00001; 
		6073: oled_colour = 16'b00001_000001_00001; 
		6074: oled_colour = 16'b00001_000001_00001; 
		6075: oled_colour = 16'b00001_000001_00001; 
		6076: oled_colour = 16'b00001_000001_00001; 
		6077: oled_colour = 16'b00001_000001_00001; 
		6078: oled_colour = 16'b00001_000001_00001; 
		6079: oled_colour = 16'b00001_000001_00001; 
		6080: oled_colour = 16'b00001_000001_00001; 
		6081: oled_colour = 16'b00001_000001_00001; 
		6082: oled_colour = 16'b00001_000001_00001; 
		6083: oled_colour = 16'b00001_000001_00001; 
		6084: oled_colour = 16'b00001_000001_00001; 
		6085: oled_colour = 16'b00001_000001_00001; 
		6086: oled_colour = 16'b00001_000001_00001; 
		6087: oled_colour = 16'b00001_000001_00001; 
		6088: oled_colour = 16'b00001_000001_00001; 
		6089: oled_colour = 16'b00001_000001_00001; 
		6090: oled_colour = 16'b00001_000001_00001; 
		6091: oled_colour = 16'b00001_000001_00001; 
		6092: oled_colour = 16'b00001_000001_00001; 
		6093: oled_colour = 16'b00001_000001_00001; 
		6094: oled_colour = 16'b00001_000001_00001; 
		6095: oled_colour = 16'b00001_000001_00001; 
		6096: oled_colour = 16'b00001_000001_00001; 
		6097: oled_colour = 16'b00001_000001_00001; 
		6098: oled_colour = 16'b00001_000001_00001; 
		6099: oled_colour = 16'b00001_000001_00001; 
		6100: oled_colour = 16'b00001_000001_00001; 
		6101: oled_colour = 16'b00001_000001_00001; 
		6102: oled_colour = 16'b00001_000001_00001; 
		6103: oled_colour = 16'b00001_000001_00001; 
		6104: oled_colour = 16'b00001_000001_00001; 
		6105: oled_colour = 16'b00001_000001_00001; 
		6106: oled_colour = 16'b00001_000001_00001; 
		6107: oled_colour = 16'b00001_000001_00001; 
		6108: oled_colour = 16'b00001_000001_00001; 
		6109: oled_colour = 16'b00001_000001_00001; 
		6110: oled_colour = 16'b00001_000001_00001; 
		6111: oled_colour = 16'b00001_000001_00001; 
		6112: oled_colour = 16'b00001_000001_00001; 
		6113: oled_colour = 16'b00001_000001_00001; 
		6114: oled_colour = 16'b00001_000001_00001; 
		6115: oled_colour = 16'b00001_000001_00001; 
		6116: oled_colour = 16'b00001_000001_00001; 
		6117: oled_colour = 16'b00001_000001_00001; 
		6118: oled_colour = 16'b00001_000001_00001; 
		6119: oled_colour = 16'b00001_000001_00001; 
		6120: oled_colour = 16'b00001_000001_00001; 
		6121: oled_colour = 16'b00001_000001_00001; 
		6122: oled_colour = 16'b00001_000001_00001; 
		6123: oled_colour = 16'b00001_000001_00001; 
		6124: oled_colour = 16'b00001_000001_00001; 
		6125: oled_colour = 16'b00001_000001_00001; 
		6126: oled_colour = 16'b00001_000001_00001; 
		6127: oled_colour = 16'b00001_000001_00001; 
		6128: oled_colour = 16'b00001_000001_00001; 
		6129: oled_colour = 16'b00001_000001_00001; 
		6130: oled_colour = 16'b00001_000001_00001; 
		6131: oled_colour = 16'b00001_000001_00001; 
		6132: oled_colour = 16'b00001_000001_00001; 
		6133: oled_colour = 16'b00001_000001_00001; 
		6134: oled_colour = 16'b00001_000001_00001; 
		6135: oled_colour = 16'b00001_000001_00001; 
		6136: oled_colour = 16'b00001_000001_00001; 
		6137: oled_colour = 16'b00001_000001_00001; 
		6138: oled_colour = 16'b00001_000001_00001; 
		6139: oled_colour = 16'b00001_000001_00001; 
		6140: oled_colour = 16'b00001_000001_00001; 
		6141: oled_colour = 16'b00001_000001_00001; 
		6142: oled_colour = 16'b00001_000001_00001; 
		6143: oled_colour = 16'b00001_000001_00001; 
		default: oled_colour = 16'b00000_000000_00000; 
	endcase
end

endmodule