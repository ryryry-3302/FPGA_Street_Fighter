module Gui_Inj3(
    input [12:0] pixel_index, 
    output reg [15:0] oled_colour 
); 

always@(pixel_index) 
begin
	case(pixel_index)
		1776: oled_colour = 16'b11110_111011_11110; 
		1777: oled_colour = 16'b11110_111010_11001; 
		1873: oled_colour = 16'b11100_110001_10000; 
		1874: oled_colour = 16'b11101_110111_01000; 
		1875: oled_colour = 16'b11110_111011_10110; 
		1876: oled_colour = 16'b11111_111110_11111; 
		1962: oled_colour = 16'b11111_111110_11111; 
		1963: oled_colour = 16'b11110_111000_11100; 
		1964: oled_colour = 16'b11011_110111_11011; 
		1965: oled_colour = 16'b10111_110010_11000; 
		1966: oled_colour = 16'b10110_110000_10110; 
		1967: oled_colour = 16'b10110_101011_10100; 
		1968: oled_colour = 16'b11010_101110_10110; 
		1969: oled_colour = 16'b11110_110100_01101; 
		1970: oled_colour = 16'b11101_110001_00111; 
		1971: oled_colour = 16'b11101_110100_00101; 
		1972: oled_colour = 16'b11101_110111_01110; 
		1973: oled_colour = 16'b11111_111100_11110; 
		2057: oled_colour = 16'b11100_110100_11010; 
		2058: oled_colour = 16'b11010_101000_10001; 
		2059: oled_colour = 16'b11100_101100_10001; 
		2060: oled_colour = 16'b10101_100000_01011; 
		2061: oled_colour = 16'b01100_100110_01100; 
		2062: oled_colour = 16'b01100_100000_01000; 
		2063: oled_colour = 16'b10010_011010_00111; 
		2064: oled_colour = 16'b11000_100011_01010; 
		2065: oled_colour = 16'b11110_110110_00111; 
		2066: oled_colour = 16'b11110_110100_01000; 
		2067: oled_colour = 16'b11101_110000_01000; 
		2068: oled_colour = 16'b11110_110100_00110; 
		2069: oled_colour = 16'b11101_110110_01000; 
		2070: oled_colour = 16'b11110_111001_11010; 
		2152: oled_colour = 16'b11101_111010_11101; 
		2153: oled_colour = 16'b11001_100100_01111; 
		2154: oled_colour = 16'b11110_110010_10010; 
		2155: oled_colour = 16'b11111_111010_11010; 
		2156: oled_colour = 16'b11011_101011_10100; 
		2157: oled_colour = 16'b01110_011011_01000; 
		2158: oled_colour = 16'b01011_011010_00111; 
		2159: oled_colour = 16'b10110_100000_01011; 
		2160: oled_colour = 16'b11001_100101_01110; 
		2161: oled_colour = 16'b11001_100101_01011; 
		2162: oled_colour = 16'b11011_101000_01110; 
		2163: oled_colour = 16'b11101_110010_10001; 
		2164: oled_colour = 16'b11101_101111_01001; 
		2165: oled_colour = 16'b11110_110010_01000; 
		2166: oled_colour = 16'b11100_101110_01010; 
		2167: oled_colour = 16'b11011_101111_10111; 
		2168: oled_colour = 16'b11111_111110_11111; 
		2248: oled_colour = 16'b10111_101101_10100; 
		2249: oled_colour = 16'b11001_100001_01100; 
		2250: oled_colour = 16'b11101_101111_10010; 
		2251: oled_colour = 16'b11101_100110_01100; 
		2252: oled_colour = 16'b10111_100010_10000; 
		2253: oled_colour = 16'b11000_100011_01110; 
		2254: oled_colour = 16'b01101_100010_01100; 
		2255: oled_colour = 16'b10000_011010_00111; 
		2256: oled_colour = 16'b10111_100010_01100; 
		2257: oled_colour = 16'b11011_101010_10001; 
		2258: oled_colour = 16'b11001_101011_10011; 
		2259: oled_colour = 16'b11001_101000_10010; 
		2260: oled_colour = 16'b11011_101110_10001; 
		2261: oled_colour = 16'b11110_110010_01100; 
		2262: oled_colour = 16'b11011_101101_01100; 
		2263: oled_colour = 16'b11001_101010_10101; 
		2344: oled_colour = 16'b01111_100011_01101; 
		2345: oled_colour = 16'b10110_011101_01010; 
		2346: oled_colour = 16'b11010_100111_01110; 
		2347: oled_colour = 16'b11110_110011_10100; 
		2348: oled_colour = 16'b11111_110010_10011; 
		2349: oled_colour = 16'b11101_101110_10000; 
		2350: oled_colour = 16'b10100_101001_01111; 
		2351: oled_colour = 16'b01101_100011_01011; 
		2352: oled_colour = 16'b10101_100000_01011; 
		2353: oled_colour = 16'b11001_101010_10010; 
		2354: oled_colour = 16'b11000_101001_10001; 
		2355: oled_colour = 16'b11010_100110_01110; 
		2356: oled_colour = 16'b11110_110001_10011; 
		2357: oled_colour = 16'b11101_110100_10111; 
		2358: oled_colour = 16'b11100_101100_10001; 
		2359: oled_colour = 16'b11100_101100_10000; 
		2360: oled_colour = 16'b11011_101111_10110; 
		2361: oled_colour = 16'b11111_111110_11111; 
		2440: oled_colour = 16'b01011_100000_01011; 
		2441: oled_colour = 16'b10001_011101_01000; 
		2442: oled_colour = 16'b11001_100000_01100; 
		2443: oled_colour = 16'b11100_101110_10100; 
		2444: oled_colour = 16'b11110_110101_10110; 
		2445: oled_colour = 16'b11110_101101_10000; 
		2446: oled_colour = 16'b11011_100110_01111; 
		2447: oled_colour = 16'b10110_101000_01111; 
		2448: oled_colour = 16'b10000_011110_01001; 
		2449: oled_colour = 16'b10001_100010_01011; 
		2450: oled_colour = 16'b01100_100011_01100; 
		2451: oled_colour = 16'b10100_011111_01100; 
		2452: oled_colour = 16'b11001_100010_01101; 
		2453: oled_colour = 16'b11001_101000_01111; 
		2454: oled_colour = 16'b11000_100011_01101; 
		2455: oled_colour = 16'b11101_110010_10100; 
		2456: oled_colour = 16'b11110_110000_10001; 
		2457: oled_colour = 16'b11010_101011_10100; 
		2536: oled_colour = 16'b10001_101010_10010; 
		2537: oled_colour = 16'b00101_011000_00100; 
		2538: oled_colour = 16'b01000_010111_00100; 
		2539: oled_colour = 16'b01100_010111_00101; 
		2540: oled_colour = 16'b10111_100100_01101; 
		2541: oled_colour = 16'b11111_110010_10011; 
		2542: oled_colour = 16'b11110_101111_10001; 
		2543: oled_colour = 16'b11111_110101_10110; 
		2544: oled_colour = 16'b11110_110101_10111; 
		2545: oled_colour = 16'b11010_101011_10000; 
		2546: oled_colour = 16'b10011_100010_01100; 
		2547: oled_colour = 16'b11011_110101_11100; 
		2548: oled_colour = 16'b11001_101100_10101; 
		2549: oled_colour = 16'b10110_011111_01010; 
		2550: oled_colour = 16'b10111_100001_01100; 
		2551: oled_colour = 16'b11000_100100_01100; 
		2552: oled_colour = 16'b11010_100101_01101; 
		2553: oled_colour = 16'b11001_100110_10001; 
		2554: oled_colour = 16'b11111_111101_11111; 
		2632: oled_colour = 16'b10111_101011_10100; 
		2633: oled_colour = 16'b01010_010100_00011; 
		2634: oled_colour = 16'b00101_010111_00011; 
		2635: oled_colour = 16'b00010_010101_00001; 
		2636: oled_colour = 16'b00110_010111_00011; 
		2637: oled_colour = 16'b10110_100110_01110; 
		2638: oled_colour = 16'b11010_101001_10001; 
		2639: oled_colour = 16'b11010_101010_10010; 
		2640: oled_colour = 16'b11000_100111_10000; 
		2641: oled_colour = 16'b11010_100101_01110; 
		2642: oled_colour = 16'b11101_101001_10000; 
		2643: oled_colour = 16'b11011_101010_10001; 
		2644: oled_colour = 16'b11011_110010_11001; 
		2645: oled_colour = 16'b11100_110110_11011; 
		2646: oled_colour = 16'b11000_100110_10001; 
		2647: oled_colour = 16'b11000_100110_10001; 
		2648: oled_colour = 16'b11010_101110_10111; 
		2649: oled_colour = 16'b11111_111110_11111; 
		2727: oled_colour = 16'b11110_111101_11111; 
		2728: oled_colour = 16'b01011_011111_01011; 
		2729: oled_colour = 16'b10010_011110_01011; 
		2730: oled_colour = 16'b11010_100111_01111; 
		2731: oled_colour = 16'b10101_011101_01010; 
		2732: oled_colour = 16'b10011_011101_01001; 
		2733: oled_colour = 16'b11001_101111_10010; 
		2734: oled_colour = 16'b10001_100001_01101; 
		2735: oled_colour = 16'b11110_111011_11110; 
		2736: oled_colour = 16'b11111_111110_11111; 
		2737: oled_colour = 16'b11010_101100_10100; 
		2738: oled_colour = 16'b10111_011111_01011; 
		2739: oled_colour = 16'b10111_100001_01011; 
		2740: oled_colour = 16'b11000_100100_01111; 
		2823: oled_colour = 16'b11100_111001_11101; 
		2824: oled_colour = 16'b01111_011010_01001; 
		2825: oled_colour = 16'b10101_100001_01101; 
		2826: oled_colour = 16'b10110_100100_01110; 
		2827: oled_colour = 16'b10100_101101_10001; 
		2828: oled_colour = 16'b10001_100000_01001; 
		2829: oled_colour = 16'b01111_100100_01100; 
		2830: oled_colour = 16'b01010_011110_00111; 
		2831: oled_colour = 16'b10000_100100_01111; 
		2834: oled_colour = 16'b11011_110000_10111; 
		2835: oled_colour = 16'b11100_110101_11010; 
		2836: oled_colour = 16'b11110_111010_11101; 
		2919: oled_colour = 16'b11110_111100_11110; 
		2920: oled_colour = 16'b01110_011011_01001; 
		2921: oled_colour = 16'b01101_100010_01100; 
		2922: oled_colour = 16'b01100_100101_01101; 
		2923: oled_colour = 16'b01011_100111_01101; 
		2924: oled_colour = 16'b10001_101101_01111; 
		2925: oled_colour = 16'b01111_100110_01101; 
		2926: oled_colour = 16'b01011_100011_01100; 
		2927: oled_colour = 16'b01100_100101_01010; 
		2928: oled_colour = 16'b10010_101011_10001; 
		2929: oled_colour = 16'b11001_110011_11001; 
		3016: oled_colour = 16'b10001_101001_10010; 
		3017: oled_colour = 16'b01001_100000_01010; 
		3018: oled_colour = 16'b01100_100101_01100; 
		3019: oled_colour = 16'b01001_011111_01001; 
		3020: oled_colour = 16'b11000_110110_10101; 
		3021: oled_colour = 16'b11000_110101_10110; 
		3022: oled_colour = 16'b01001_011100_00111; 
		3023: oled_colour = 16'b01111_011110_00111; 
		3024: oled_colour = 16'b11101_110001_10010; 
		3025: oled_colour = 16'b10110_101100_10011; 
		3026: oled_colour = 16'b11011_110111_11100; 
		3112: oled_colour = 16'b11110_111100_11111; 
		3113: oled_colour = 16'b01100_100001_01100; 
		3114: oled_colour = 16'b10000_101011_10000; 
		3115: oled_colour = 16'b10010_101100_10010; 
		3116: oled_colour = 16'b11000_101110_10010; 
		3117: oled_colour = 16'b11111_111101_11101; 
		3118: oled_colour = 16'b10111_110010_10110; 
		3119: oled_colour = 16'b10011_101100_01111; 
		3120: oled_colour = 16'b11011_111000_10101; 
		3121: oled_colour = 16'b11111_111111_11100; 
		3122: oled_colour = 16'b10101_101110_10010; 
		3123: oled_colour = 16'b10010_101001_10011; 
		3124: oled_colour = 16'b11111_111110_11111; 
		3209: oled_colour = 16'b10101_101110_10101; 
		3210: oled_colour = 16'b10010_100010_01101; 
		3211: oled_colour = 16'b11000_110001_10100; 
		3213: oled_colour = 16'b11110_111100_11101; 
		3214: oled_colour = 16'b11101_111011_11010; 
		3215: oled_colour = 16'b01110_101001_01110; 
		3216: oled_colour = 16'b10011_101111_10001; 
		3217: oled_colour = 16'b11110_111001_10111; 
		3218: oled_colour = 16'b11110_111111_11010; 
		3219: oled_colour = 16'b10011_110000_10001; 
		3220: oled_colour = 16'b10001_101000_10001; 
		3305: oled_colour = 16'b11001_110100_11010; 
		3306: oled_colour = 16'b01110_011010_01001; 
		3307: oled_colour = 16'b11011_110101_11001; 
		3308: oled_colour = 16'b10111_110100_10111; 
		3309: oled_colour = 16'b11000_110100_10010; 
		3310: oled_colour = 16'b11111_111001_11000; 
		3311: oled_colour = 16'b10010_101011_01111; 
		3312: oled_colour = 16'b01101_100011_01101; 
		3313: oled_colour = 16'b11000_110111_11001; 
		3314: oled_colour = 16'b11000_111010_10101; 
		3315: oled_colour = 16'b11110_111111_11001; 
		3316: oled_colour = 16'b10001_101110_10001; 
		3317: oled_colour = 16'b11011_110111_11100; 
		3402: oled_colour = 16'b10110_110000_10111; 
		3403: oled_colour = 16'b01101_100010_01100; 
		3404: oled_colour = 16'b01011_011111_01010; 
		3405: oled_colour = 16'b10101_110110_10010; 
		3406: oled_colour = 16'b11111_111111_11100; 
		3407: oled_colour = 16'b11010_111011_11001; 
		3408: oled_colour = 16'b01010_100001_01010; 
		3409: oled_colour = 16'b01110_100001_01011; 
		3410: oled_colour = 16'b10110_110010_10010; 
		3411: oled_colour = 16'b11011_111001_10100; 
		3412: oled_colour = 16'b10110_101110_10000; 
		3413: oled_colour = 16'b11001_110000_11000; 
		3497: oled_colour = 16'b11011_111000_11100; 
		3498: oled_colour = 16'b01011_011110_01010; 
		3499: oled_colour = 16'b01100_010111_00110; 
		3500: oled_colour = 16'b01101_010111_00101; 
		3501: oled_colour = 16'b10100_101101_01110; 
		3502: oled_colour = 16'b11110_111111_11011; 
		3503: oled_colour = 16'b11001_111010_11000; 
		3504: oled_colour = 16'b01000_011101_00111; 
		3505: oled_colour = 16'b10010_011101_01011; 
		3506: oled_colour = 16'b11101_101010_10000; 
		3507: oled_colour = 16'b11110_110000_10010; 
		3508: oled_colour = 16'b11010_100101_01110; 
		3509: oled_colour = 16'b11010_110000_11000; 
		3592: oled_colour = 16'b11110_111100_11110; 
		3593: oled_colour = 16'b01100_010101_00101; 
		3594: oled_colour = 16'b10001_101000_10001; 
		3595: oled_colour = 16'b11100_111000_11001; 
		3596: oled_colour = 16'b11010_101101_10000; 
		3597: oled_colour = 16'b11110_110010_10011; 
		3598: oled_colour = 16'b11011_110100_10101; 
		3599: oled_colour = 16'b10000_101000_01110; 
		3600: oled_colour = 16'b01010_011001_00111; 
		3601: oled_colour = 16'b01010_011110_01010; 
		3602: oled_colour = 16'b10100_110110_10100; 
		3603: oled_colour = 16'b11110_111111_11000; 
		3604: oled_colour = 16'b10101_110001_10010; 
		3605: oled_colour = 16'b10111_110010_11000; 
		3688: oled_colour = 16'b11010_110101_11010; 
		3689: oled_colour = 16'b00110_001110_00001; 
		3690: oled_colour = 16'b10100_101100_10000; 
		3691: oled_colour = 16'b11111_111111_11101; 
		3692: oled_colour = 16'b11100_111011_11000; 
		3693: oled_colour = 16'b10011_101000_01110; 
		3694: oled_colour = 16'b10100_100001_01110; 
		3695: oled_colour = 16'b11100_110110_11011; 
		3696: oled_colour = 16'b11100_110101_11010; 
		3697: oled_colour = 16'b01001_010001_00010; 
		3698: oled_colour = 16'b01110_100100_01011; 
		3699: oled_colour = 16'b10111_111001_10100; 
		3700: oled_colour = 16'b01110_101010_01110; 
		3701: oled_colour = 16'b10110_110000_10111; 
		3784: oled_colour = 16'b10110_100010_01111; 
		3785: oled_colour = 16'b10000_011101_01000; 
		3786: oled_colour = 16'b01010_100000_01000; 
		3787: oled_colour = 16'b10010_101101_10000; 
		3788: oled_colour = 16'b01110_100111_01110; 
		3789: oled_colour = 16'b10101_101111_10110; 
		3793: oled_colour = 16'b10000_100100_01110; 
		3794: oled_colour = 16'b01001_010011_00010; 
		3795: oled_colour = 16'b01100_011101_01001; 
		3796: oled_colour = 16'b01011_011000_00110; 
		3797: oled_colour = 16'b11011_110111_11011; 
		3879: oled_colour = 16'b10100_100011_01111; 
		3880: oled_colour = 16'b01101_010000_00001; 
		3881: oled_colour = 16'b10101_011101_01010; 
		3882: oled_colour = 16'b01111_010110_00101; 
		3883: oled_colour = 16'b01111_100000_01100; 
		3884: oled_colour = 16'b11110_111011_11110; 
		3889: oled_colour = 16'b11101_111001_11101; 
		3890: oled_colour = 16'b10011_011010_01001; 
		3891: oled_colour = 16'b10100_011010_01000; 
		3892: oled_colour = 16'b10011_011010_01000; 
		3893: oled_colour = 16'b11111_111100_11110; 
		3974: oled_colour = 16'b11010_101101_10110; 
		3975: oled_colour = 16'b10011_011001_00111; 
		3976: oled_colour = 16'b01011_010000_00001; 
		3977: oled_colour = 16'b01111_010100_00100; 
		3978: oled_colour = 16'b10111_100101_10000; 
		3985: oled_colour = 16'b11100_111000_11100; 
		3986: oled_colour = 16'b01011_001111_00001; 
		3987: oled_colour = 16'b01101_010001_00010; 
		3988: oled_colour = 16'b10010_011001_01000; 
		3989: oled_colour = 16'b11111_111100_11110; 
		4070: oled_colour = 16'b11011_101100_10011; 
		4071: oled_colour = 16'b10010_010111_00101; 
		4072: oled_colour = 16'b01100_010001_00010; 
		4073: oled_colour = 16'b10101_011110_01011; 
		4074: oled_colour = 16'b11101_111001_11110; 
		4081: oled_colour = 16'b11001_101011_10100; 
		4082: oled_colour = 16'b10000_010100_00100; 
		4083: oled_colour = 16'b01101_010010_00010; 
		4084: oled_colour = 16'b10010_011001_01000; 
		4085: oled_colour = 16'b11100_110110_11011; 
		4167: oled_colour = 16'b11001_101101_10101; 
		4168: oled_colour = 16'b01110_010011_00100; 
		4169: oled_colour = 16'b10110_011110_01010; 
		4170: oled_colour = 16'b11000_100100_01110; 
		4171: oled_colour = 16'b11100_110100_11010; 
		4177: oled_colour = 16'b11010_101010_10011; 
		4178: oled_colour = 16'b10101_011011_01001; 
		4179: oled_colour = 16'b01011_001110_00001; 
		4180: oled_colour = 16'b01111_010011_00100; 
		4181: oled_colour = 16'b10101_011111_01100; 
		4182: oled_colour = 16'b11011_101110_10110; 
		4183: oled_colour = 16'b11111_111100_11110; 
		4264: oled_colour = 16'b11100_110100_11010; 
		4265: oled_colour = 16'b11010_101001_10010; 
		4266: oled_colour = 16'b11010_101100_10100; 
		4267: oled_colour = 16'b11010_101110_10111; 
		4273: oled_colour = 16'b11111_111100_11110; 
		4274: oled_colour = 16'b11101_111000_11100; 
		4275: oled_colour = 16'b11000_101100_10101; 
		4276: oled_colour = 16'b10100_011101_01100; 
		4277: oled_colour = 16'b11000_100100_01111; 
		4278: oled_colour = 16'b11000_100011_01110; 
		4279: oled_colour = 16'b11011_110010_11001; 
		4373: oled_colour = 16'b11111_111101_11111; 
		4374: oled_colour = 16'b11111_111110_11111; 
		default: oled_colour = 16'b00000_000000_00000; 
	endcase
end

endmodule