
module HealthManagement (input clk, output reg [5:0]health_1, output reg [5:0] health_2)


endmodule
```
